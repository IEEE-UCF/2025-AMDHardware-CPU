// System Control Coprocessor (CP0)
// Handles system-level operations like CSR access, exceptions, and privileged instructions

module coprocessor_cp0 #(
    parameter ADDR_WIDTH = 64,
    parameter DATA_WIDTH = 64,
    parameter INST_WIDTH = 32
)(
    input  logic                    clk,
    input  logic                    rst_n,
    
    // Coprocessor Interface
    input  logic                    cp_enable,
    input  logic [INST_WIDTH-1:0]  cp_instruction,
    input  logic [DATA_WIDTH-1:0]  cp_data_in,
    output logic [DATA_WIDTH-1:0]  cp_data_out,
    output logic                    cp_ready,
    output logic                    cp_exception,
    
    // System Interface
    input  logic                    interrupt_pending,
    input  logic [DATA_WIDTH-1:0]  pc_current,
    output logic                    trap_enable,
    output logic [DATA_WIDTH-1:0]  trap_vector,
    output logic                    privilege_mode,  // 0=user, 1=supervisor
    
    // Debug Interface
    output logic                    debug_mode,
    output logic [DATA_WIDTH-1:0]  debug_pc
);

    // CSR (Control and Status Register) definitions
    typedef enum logic [11:0] {
        CSR_MSTATUS   = 12'h300,  // Machine status
        CSR_MISA      = 12'h301,  // Machine ISA
        CSR_MIE       = 12'h304,  // Machine interrupt enable
        CSR_MTVEC     = 12'h305,  // Machine trap vector
        CSR_MSCRATCH  = 12'h340,  // Machine scratch
        CSR_MEPC      = 12'h341,  // Machine exception PC
        CSR_MCAUSE    = 12'h342,  // Machine cause
        CSR_MTVAL     = 12'h343,  // Machine trap value
        CSR_MIP       = 12'h344,  // Machine interrupt pending
        CSR_CYCLE     = 12'hC00,  // Cycle counter
        CSR_INSTRET   = 12'hC02   // Instructions retired
    } csr_addr_t;

    // CSR registers
    logic [DATA_WIDTH-1:0] csr_mstatus;
    logic [DATA_WIDTH-1:0] csr_misa;
    logic [DATA_WIDTH-1:0] csr_mie;
    logic [DATA_WIDTH-1:0] csr_mtvec;
    logic [DATA_WIDTH-1:0] csr_mscratch;
    logic [DATA_WIDTH-1:0] csr_mepc;
    logic [DATA_WIDTH-1:0] csr_mcause;
    logic [DATA_WIDTH-1:0] csr_mtval;
    logic [DATA_WIDTH-1:0] csr_mip;
    logic [DATA_WIDTH-1:0] csr_cycle;
    logic [DATA_WIDTH-1:0] csr_instret;
    
    // Instruction decode
    logic [6:0]  opcode;
    logic [2:0]  funct3;
    logic [11:0] csr_addr;
    logic [4:0]  rs1;
    logic [4:0]  rd;
    logic [4:0]  zimm;
    
    assign opcode = cp_instruction[6:0];
    assign funct3 = cp_instruction[14:12];
    assign csr_addr = cp_instruction[31:20];
    assign rs1 = cp_instruction[19:15];
    assign rd = cp_instruction[11:7];
    assign zimm = cp_instruction[19:15]; // Zero-extended immediate for CSRR*I
    
    // CSR operation types
    typedef enum logic [2:0] {
        CSR_RW   = 3'b001,  // CSRRW
        CSR_RS   = 3'b010,  // CSRRS
        CSR_RC   = 3'b011,  // CSRRC
        CSR_RWI  = 3'b101,  // CSRRWI
        CSR_RSI  = 3'b110,  // CSRRSI
        CSR_RCI  = 3'b111   // CSRRCI
    } csr_op_t;
    
    // Internal signals
    logic csr_write_enable;
    logic [DATA_WIDTH-1:0] csr_write_data;
    logic [DATA_WIDTH-1:0] csr_read_data;
    logic csr_valid;
    logic is_csr_instruction;
    logic is_immediate_op;
    
    // Detect CSR instructions (SYSTEM opcode)
    assign is_csr_instruction = cp_enable && (opcode == 7'b1110011) && (funct3 != 3'b000);
    assign is_immediate_op = funct3[2]; // Bit 2 indicates immediate operation
    assign csr_valid = is_csr_instruction;
    
    // CSR read logic
    always_comb begin
        csr_read_data = '0;
        case (csr_addr)
            CSR_MSTATUS:  csr_read_data = csr_mstatus;
            CSR_MISA:     csr_read_data = csr_misa;
            CSR_MIE:      csr_read_data = csr_mie;
            CSR_MTVEC:    csr_read_data = csr_mtvec;
            CSR_MSCRATCH: csr_read_data = csr_mscratch;
            CSR_MEPC:     csr_read_data = csr_mepc;
            CSR_MCAUSE:   csr_read_data = csr_mcause;
            CSR_MTVAL:    csr_read_data = csr_mtval;
            CSR_MIP:      csr_read_data = csr_mip;
            CSR_CYCLE:    csr_read_data = csr_cycle;
            CSR_INSTRET:  csr_read_data = csr_instret;
            default:      csr_read_data = '0;
        endcase
    end
    
    // CSR write data calculation
    always_comb begin
        csr_write_enable = 1'b0;
        csr_write_data = '0;
        
        if (csr_valid) begin
            case (funct3)
                CSR_RW, CSR_RWI: begin
                    csr_write_enable = 1'b1;
                    csr_write_data = is_immediate_op ? {{(DATA_WIDTH-5){1'b0}}, zimm} : cp_data_in;
                end
                CSR_RS, CSR_RSI: begin
                    csr_write_enable = (is_immediate_op ? (zimm != 0) : (rs1 != 0));
                    csr_write_data = csr_read_data | (is_immediate_op ? {{(DATA_WIDTH-5){1'b0}}, zimm} : cp_data_in);
                end
                CSR_RC, CSR_RCI: begin
                    csr_write_enable = (is_immediate_op ? (zimm != 0) : (rs1 != 0));
                    csr_write_data = csr_read_data & ~(is_immediate_op ? {{(DATA_WIDTH-5){1'b0}}, zimm} : cp_data_in);
                end
                default: begin
                    csr_write_enable = 1'b0;
                    csr_write_data = '0;
                end
            endcase
        end
    end
    
    // CSR register updates
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            csr_mstatus <= '0;
            csr_misa <= 64'h8000000000141101; // RV64I with some extensions
            csr_mie <= '0;
            csr_mtvec <= '0;
            csr_mscratch <= '0;
            csr_mepc <= '0;
            csr_mcause <= '0;
            csr_mtval <= '0;
            csr_mip <= '0;
            csr_cycle <= '0;
            csr_instret <= '0;
        end else begin
            // Update cycle and instruction counters
            csr_cycle <= csr_cycle + 1;
            if (cp_enable) begin
                csr_instret <= csr_instret + 1;
            end
            
            // Handle interrupt pending
            csr_mip[7] <= interrupt_pending; // Machine timer interrupt
            
            // CSR writes
            if (csr_write_enable) begin
                case (csr_addr)
                    CSR_MSTATUS:  csr_mstatus <= csr_write_data;
                    CSR_MIE:      csr_mie <= csr_write_data;
                    CSR_MTVEC:    csr_mtvec <= csr_write_data;
                    CSR_MSCRATCH: csr_mscratch <= csr_write_data;
                    CSR_MEPC:     csr_mepc <= csr_write_data;
                    CSR_MCAUSE:   csr_mcause <= csr_write_data;
                    CSR_MTVAL:    csr_mtval <= csr_write_data;
                    default: ; // Read-only or invalid CSR
                endcase
            end
        end
    end
    
    // Output assignments
    assign cp_data_out = csr_read_data;
    assign cp_ready = 1'b1; // CSR operations complete in one cycle
    assign cp_exception = csr_valid && (csr_addr == 12'h000); // Invalid CSR address
    
    // System control outputs
    assign trap_enable = interrupt_pending && csr_mie[7] && csr_mstatus[3]; // Machine interrupt enable
    assign trap_vector = csr_mtvec;
    assign privilege_mode = csr_mstatus[3]; // Machine mode
    assign debug_mode = 1'b0; // Not implemented in this basic version
    assign debug_pc = pc_current;

endmodule

// Floating Point Coprocessor (CP1)
// Handles floating point arithmetic operations

module coprocessor_cp1 #(
    parameter ADDR_WIDTH = 64,
    parameter DATA_WIDTH = 64,
    parameter INST_WIDTH = 32,
    parameter FP_REG_NUM = 32
)(
    input  logic                    clk,
    input  logic                    rst_n,
    
    // Coprocessor Interface
    input  logic                    cp_enable,
    input  logic [INST_WIDTH-1:0]  cp_instruction,
    input  logic [DATA_WIDTH-1:0]  cp_data_in,
    output logic [DATA_WIDTH-1:0]  cp_data_out,
    output logic                    cp_ready,
    output logic                    cp_exception,
    
    // Floating Point Register File Interface
    output logic                    fp_reg_write,
    output logic [4:0]              fp_reg_waddr,
    output logic [DATA_WIDTH-1:0]   fp_reg_wdata,
    output logic [4:0]              fp_reg_raddr1,
    output logic [4:0]              fp_reg_raddr2,
    input  logic [DATA_WIDTH-1:0]   fp_reg_rdata1,
    input  logic [DATA_WIDTH-1:0]   fp_reg_rdata2,
    
    // Status flags
    output logic                    fp_invalid,
    output logic                    fp_divide_by_zero,
    output logic                    fp_overflow,
    output logic                    fp_underflow,
    output logic                    fp_inexact
);

    // Instruction decode
    logic [6:0]  opcode;
    logic [4:0]  rd, rs1, rs2;
    logic [2:0]  funct3;
    logic [6:0]  funct7;
    logic [4:0]  rs3;
    logic [1:0]  fmt;        // Format: 00=S(32-bit), 01=D(64-bit)
    logic [2:0]  rm;         // Rounding mode
    
    assign opcode = cp_instruction[6:0];
    assign rd = cp_instruction[11:7];
    assign funct3 = cp_instruction[14:12];
    assign rs1 = cp_instruction[19:15];
    assign rs2 = cp_instruction[24:20];
    assign funct7 = cp_instruction[31:25];
    assign rs3 = cp_instruction[31:27];
    assign fmt = cp_instruction[26:25];
    assign rm = cp_instruction[14:12];
    
    // FP operation types
    typedef enum logic [6:0] {
        FP_LOAD     = 7'b0000111,  // FLW, FLD
        FP_STORE    = 7'b0100111,  // FSW, FSD
        FP_MADD     = 7'b1000011,  // FMADD
        FP_MSUB     = 7'b1000111,  // FMSUB
        FP_NMSUB    = 7'b1001011,  // FNMSUB
        FP_NMADD    = 7'b1001111,  // FNMADD
        FP_OP       = 7'b1010011   // FP arithmetic
    } fp_opcode_t;
    
    // FP arithmetic function codes
    typedef enum logic [6:0] {
        FP_ADD      = 7'b0000000,  // FADD
        FP_SUB      = 7'b0000100,  // FSUB
        FP_MUL      = 7'b0001000,  // FMUL
        FP_DIV      = 7'b0001100,  // FDIV
        FP_SQRT     = 7'b0101100,  // FSQRT
        FP_SGNJ     = 7'b0010000,  // FSGNJ, FSGNJN, FSGNJX
        FP_MINMAX   = 7'b0010100,  // FMIN, FMAX
        FP_CVT_W    = 7'b1100000,  // FCVT.W.S/D
        FP_CVT_WU   = 7'b1100001,  // FCVT.WU.S/D
        FP_CVT_L    = 7'b1100010,  // FCVT.L.S/D
        FP_CVT_LU   = 7'b1100011,  // FCVT.LU.S/D
        FP_CVT_S    = 7'b1101000,  // FCVT.S.W/WU/L/LU
        FP_CVT_D    = 7'b1101001,  // FCVT.D.W/WU/L/LU
        FP_CVT_SD   = 7'b0100000,  // FCVT.S.D, FCVT.D.S
        FP_CMP      = 7'b1010000,  // FEQ, FLT, FLE
        FP_CLASS    = 7'b1110000,  // FCLASS
        FP_MV       = 7'b1111000   // FMV.X.W/D, FMV.W/D.X
    } fp_funct7_t;
    
    // Pipeline stages
    typedef enum logic [2:0] {
        FP_IDLE,
        FP_DECODE,
        FP_EXECUTE,
        FP_COMPLETE
    } fp_state_t;
    
    fp_state_t current_state, next_state;
    
    // Internal registers
    logic [DATA_WIDTH-1:0] operand_a, operand_b, operand_c;
    logic [DATA_WIDTH-1:0] result;
    logic result_valid;
    logic [4:0] operation_cycles;
    logic [4:0] cycle_counter;
    
    // Floating point flags
    logic fp_flags_invalid, fp_flags_div_zero, fp_flags_overflow;
    logic fp_flags_underflow, fp_flags_inexact;
    
    // Detect FP instructions
    logic is_fp_instruction;
    assign is_fp_instruction = cp_enable && (
        opcode == FP_LOAD || opcode == FP_STORE || opcode == FP_MADD ||
        opcode == FP_MSUB || opcode == FP_NMSUB || opcode == FP_NMADD ||
        opcode == FP_OP
    );
    
    // State machine
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            current_state <= FP_IDLE;
            cycle_counter <= '0;
        end else begin
            current_state <= next_state;
            if (current_state == FP_EXECUTE) begin
                cycle_counter <= cycle_counter + 1;
            end else begin
                cycle_counter <= '0;
            end
        end
    end
    
    // Next state logic
    always_comb begin
        next_state = current_state;
        case (current_state)
            FP_IDLE: begin
                if (is_fp_instruction)
                    next_state = FP_DECODE;
            end
            FP_DECODE: begin
                next_state = FP_EXECUTE;
            end
            FP_EXECUTE: begin
                if (cycle_counter >= operation_cycles)
                    next_state = FP_COMPLETE;
            end
            FP_COMPLETE: begin
                next_state = FP_IDLE;
            end
        endcase
    end
    
    // Operation cycle determination
    always_comb begin
        operation_cycles = 5'd1; // Default single cycle
        if (opcode == FP_OP) begin
            case (funct7)
                FP_ADD, FP_SUB:     operation_cycles = 5'd3;
                FP_MUL:             operation_cycles = 5'd4;
                FP_DIV:             operation_cycles = 5'd16;
                FP_SQRT:            operation_cycles = 5'd20;
                FP_CVT_W, FP_CVT_WU,
                FP_CVT_L, FP_CVT_LU,
                FP_CVT_S, FP_CVT_D,
                FP_CVT_SD:          operation_cycles = 5'd2;
                default:            operation_cycles = 5'd1;
            endcase
        end
    end
    
    // Operand selection
    always_comb begin
        operand_a = fp_reg_rdata1;
        operand_b = fp_reg_rdata2;
        operand_c = '0; // For fused multiply-add operations
        
        // Special cases for immediate operations or CPU data
        if (opcode == FP_LOAD || (opcode == FP_OP && funct7 == FP_MV && rs2[0])) begin
            operand_a = cp_data_in;
        end
    end
    
    // Simplified FP execution (placeholder for actual FP units)
    always_comb begin
        result = '0;
        fp_flags_invalid = 1'b0;
        fp_flags_div_zero = 1'b0;
        fp_flags_overflow = 1'b0;
        fp_flags_underflow = 1'b0;
        fp_flags_inexact = 1'b0;
        
        if (current_state == FP_EXECUTE || current_state == FP_COMPLETE) begin
            case (opcode)
                FP_LOAD: begin
                    result = operand_a;
                end
                FP_STORE: begin
                    result = operand_a;
                end
                FP_OP: begin
                    case (funct7)
                        FP_ADD: begin
                            // Simplified: just pass through for now
                            result = operand_a;
                        end
                        FP_SUB: begin
                            result = operand_a;
                        end
                        FP_MUL: begin
                            result = operand_a;
                        end
                        FP_DIV: begin
                            result = operand_a;
                            // Check for divide by zero
                            if (operand_b == '0) begin
                                fp_flags_div_zero = 1'b1;
                            end
                        end
                        FP_MV: begin
                            if (rs2[0]) // FMV.W/D.X
                                result = operand_a;
                            else        // FMV.X.W/D
                                result = operand_a;
                        end
                        FP_CMP: begin
                            // Comparison result (0 or 1)
                            case (funct3)
                                3'b010: result = (operand_a == operand_b) ? 1 : 0; // FEQ
                                3'b001: result = (operand_a < operand_b) ? 1 : 0;  // FLT
                                3'b000: result = (operand_a <= operand_b) ? 1 : 0; // FLE
                                default: result = '0;
                            endcase
                        end
                        default: begin
                            result = operand_a;
                        end
                    endcase
                end
                default: begin
                    result = '0;
                end
            endcase
        end
    end
    
    // Register file control
    assign fp_reg_raddr1 = rs1;
    assign fp_reg_raddr2 = rs2;
    assign fp_reg_write = (current_state == FP_COMPLETE) && 
                         (opcode != FP_STORE) && (rd != 5'b00000);
    assign fp_reg_waddr = rd;
    assign fp_reg_wdata = result;
    
    // Output assignments
    assign cp_data_out = result;
    assign cp_ready = (current_state == FP_COMPLETE) || 
                     (current_state == FP_IDLE && !is_fp_instruction);
    assign cp_exception = fp_flags_invalid || fp_flags_div_zero;
    
    // Status flags
    assign fp_invalid = fp_flags_invalid;
    assign fp_divide_by_zero = fp_flags_div_zero;
    assign fp_overflow = fp_flags_overflow;
    assign fp_underflow = fp_flags_underflow;
    assign fp_inexact = fp_flags_inexact;

endmodule

// Memory Management Coprocessor (CP2)
// Handles virtual memory, TLB, and cache control operations

module coprocessor_cp2 #(
    parameter ADDR_WIDTH = 64,
    parameter DATA_WIDTH = 64,
    parameter INST_WIDTH = 32,
    parameter TLB_ENTRIES = 64,
    parameter PAGE_SIZE = 4096
)(
    input  logic                    clk,
    input  logic                    rst_n,
    
    // Coprocessor Interface
    input  logic                    cp_enable,
    input  logic [INST_WIDTH-1:0]  cp_instruction,
    input  logic [DATA_WIDTH-1:0]  cp_data_in,
    output logic [DATA_WIDTH-1:0]  cp_data_out,
    output logic                    cp_ready,
    output logic                    cp_exception,
    
    // Memory Management Interface
    input  logic [ADDR_WIDTH-1:0]  virtual_addr,
    output logic [ADDR_WIDTH-1:0]  physical_addr,
    output logic                    translation_valid,
    output logic                    page_fault,
    
    // Cache Control Interface
    output logic                    cache_flush,
    output logic                    cache_invalidate,
    output logic [ADDR_WIDTH-1:0]  cache_addr,
    
    // System Interface
    input  logic [DATA_WIDTH-1:0]  page_table_base,
    input  logic                    vm_enable,
    output logic                    tlb_miss,
    output logic                    protection_fault
);

    // TLB Entry arrays (replacing struct due to iverilog limitations)
    logic [TLB_ENTRIES-1:0]             tlb_valid;
    logic [TLB_ENTRIES-1:0]             tlb_global;
    logic [19:0]                        tlb_vpn [TLB_ENTRIES-1:0];
    logic [43:0]                        tlb_ppn [TLB_ENTRIES-1:0];
    logic [1:0]                         tlb_privilege [TLB_ENTRIES-1:0];
    logic [TLB_ENTRIES-1:0]             tlb_readable;
    logic [TLB_ENTRIES-1:0]             tlb_writable;
    logic [TLB_ENTRIES-1:0]             tlb_executable;
    logic [TLB_ENTRIES-1:0]             tlb_accessed;
    logic [TLB_ENTRIES-1:0]             tlb_dirty;
    logic [$clog2(TLB_ENTRIES)-1:0] tlb_index;
    
    // Instruction decode
    logic [6:0]  opcode;
    logic [2:0]  funct3;
    logic [11:0] funct12;
    logic [4:0]  rs1, rs2, rd;
    
    assign opcode = cp_instruction[6:0];
    assign funct3 = cp_instruction[14:12];
    assign funct12 = cp_instruction[31:20];
    assign rs1 = cp_instruction[19:15];
    assign rs2 = cp_instruction[24:20];
    assign rd = cp_instruction[11:7];
    
    // Memory management operations
    typedef enum logic [11:0] {
        MM_SFENCE_VMA   = 12'h120,  // Supervisor fence virtual memory
        MM_SFENCE_W_INVAL = 12'h180, // Supervisor fence with invalidate
        MM_HFENCE_VVMA  = 12'h220,  // Hypervisor fence virtual memory
        MM_HFENCE_GVMA  = 12'h620,  // Hypervisor fence guest virtual memory
        MM_FLUSH_CACHE  = 12'h001,  // Custom: flush cache
        MM_INVAL_CACHE  = 12'h002,  // Custom: invalidate cache
        MM_LOAD_TLB     = 12'h003,  // Custom: load TLB entry
        MM_FLUSH_TLB    = 12'h004   // Custom: flush TLB
    } mm_funct12_t;
    
    // Internal signals
    logic is_mm_instruction;
    logic tlb_hit;
    logic [$clog2(TLB_ENTRIES)-1:0] tlb_hit_index;
    logic [19:0] lookup_vpn;
    logic [43:0] lookup_ppn;
    logic mm_operation_valid;
    logic operation_complete;
    
    // Detect memory management instructions
    assign is_mm_instruction = cp_enable && (opcode == 7'b1110011) && (funct3 == 3'b000);
    
    // Virtual to physical address translation
    assign lookup_vpn = virtual_addr[31:12]; // Assuming 32-bit virtual addresses for simplicity
    
    // TLB lookup logic
    always_comb begin
        tlb_hit = 1'b0;
        tlb_hit_index = '0;
        lookup_ppn = '0;
        
        for (int i = 0; i < TLB_ENTRIES; i++) begin
            if (tlb_valid[i] && (tlb_vpn[i] == lookup_vpn)) begin
                tlb_hit = 1'b1;
                tlb_hit_index = i[$clog2(TLB_ENTRIES)-1:0];
                lookup_ppn = tlb_ppn[i];
                i = TLB_ENTRIES; // Exit loop
            end
        end
    end
    
    // Address translation
    assign physical_addr = vm_enable ? 
                          (tlb_hit ? {lookup_ppn, virtual_addr[11:0]} : virtual_addr) :
                          virtual_addr;
    assign translation_valid = !vm_enable || tlb_hit;
    assign page_fault = vm_enable && !tlb_hit;
    assign tlb_miss = vm_enable && !tlb_hit;
    
    // Protection checking
    always_comb begin
        protection_fault = 1'b0;
        if (vm_enable && tlb_hit) begin
            // Check access permissions based on operation type
            // This is simplified - real implementation would check current privilege level
            if (!tlb_writable[tlb_hit_index]) begin
                protection_fault = 1'b1; // Would need to know if this is a write operation
            end
        end
    end
    
    // TLB management operations
    logic tlb_flush_all;
    logic tlb_flush_entry;
    logic tlb_load_entry;
    logic [TLB_ENTRIES-1:0] tlb_replacement_policy;
    logic [$clog2(TLB_ENTRIES)-1:0] tlb_replace_index;
    
    // Simple replacement policy (round-robin)
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            tlb_replace_index <= '0;
        end else if (tlb_load_entry) begin
            tlb_replace_index <= tlb_replace_index + 1;
        end
    end
    
    // Memory management operation execution
    always_comb begin
        tlb_flush_all = 1'b0;
        tlb_flush_entry = 1'b0;
        tlb_load_entry = 1'b0;
        cache_flush = 1'b0;
        cache_invalidate = 1'b0;
        cache_addr = virtual_addr;
        operation_complete = 1'b1; // Most operations complete immediately
        
        if (is_mm_instruction) begin
            case (funct12)
                MM_SFENCE_VMA: begin
                    if (rs1 == 5'b00000 && rs2 == 5'b00000) begin
                        tlb_flush_all = 1'b1;
                    end else begin
                        tlb_flush_entry = 1'b1;
                    end
                end
                MM_FLUSH_CACHE: begin
                    cache_flush = 1'b1;
                end
                MM_INVAL_CACHE: begin
                    cache_invalidate = 1'b1;
                end
                MM_LOAD_TLB: begin
                    tlb_load_entry = 1'b1;
                end
                MM_FLUSH_TLB: begin
                    tlb_flush_all = 1'b1;
                end
                default: begin
                    // Unknown operation
                end
            endcase
        end
    end
    
    // TLB updates
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            // Initialize TLB - all entries invalid
            for (int i = 0; i < TLB_ENTRIES; i++) begin
                tlb_valid[i] <= 1'b0;
                tlb_global[i] <= 1'b0;
                tlb_vpn[i] <= '0;
                tlb_ppn[i] <= '0;
                tlb_privilege[i] <= 2'b00;
                tlb_readable[i] <= 1'b0;
                tlb_writable[i] <= 1'b0;
                tlb_executable[i] <= 1'b0;
                tlb_accessed[i] <= 1'b0;
                tlb_dirty[i] <= 1'b0;
            end
        end else begin
            // Handle TLB operations
            if (tlb_flush_all) begin
                for (int i = 0; i < TLB_ENTRIES; i++) begin
                    tlb_valid[i] <= 1'b0;
                end
            end else if (tlb_flush_entry) begin
                // Flush specific entry based on rs1 (VPN) and rs2 (ASID)
                for (int i = 0; i < TLB_ENTRIES; i++) begin
                    if (tlb_vpn[i] == cp_data_in[19:0]) begin
                        tlb_valid[i] <= 1'b0;
                    end
                end
            end else if (tlb_load_entry) begin
                // Load new TLB entry from cp_data_in
                // Format: {valid, global, vpn[19:0], ppn[43:0], flags}
                tlb_valid[tlb_replace_index] <= cp_data_in[63];
                tlb_global[tlb_replace_index] <= cp_data_in[62];
                tlb_vpn[tlb_replace_index] <= cp_data_in[61:42];
                tlb_ppn[tlb_replace_index] <= cp_data_in[41:0]; // Simplified
                tlb_readable[tlb_replace_index] <= 1'b1;
                tlb_writable[tlb_replace_index] <= 1'b1;
                tlb_executable[tlb_replace_index] <= 1'b1;
                tlb_privilege[tlb_replace_index] <= 2'b01; // Supervisor
            end
            
            // Update accessed/dirty bits on TLB hit
            if (tlb_hit && vm_enable) begin
                tlb_accessed[tlb_hit_index] <= 1'b1;
                // tlb_dirty[tlb_hit_index] <= write_access; // Would need write signal
            end
        end
    end
    
    // Output assignments
    assign cp_data_out = {lookup_ppn, virtual_addr[11:0]}; // Return physical address
    assign cp_ready = operation_complete;
    assign cp_exception = is_mm_instruction && (funct12 > MM_FLUSH_TLB); // Invalid operation

endmodule

// Debug Coprocessor (CP3)
// Handles debugging, performance monitoring, and trace functionality

module coprocessor_cp3 #(
    parameter ADDR_WIDTH = 64,
    parameter DATA_WIDTH = 64,
    parameter INST_WIDTH = 32,
    parameter NUM_BREAKPOINTS = 8,
    parameter NUM_WATCHPOINTS = 4,
    parameter TRACE_BUFFER_SIZE = 256
)(
    input  logic                    clk,
    input  logic                    rst_n,
    
    // Coprocessor Interface
    input  logic                    cp_enable,
    input  logic [INST_WIDTH-1:0]  cp_instruction,
    input  logic [DATA_WIDTH-1:0]  cp_data_in,
    output logic [DATA_WIDTH-1:0]  cp_data_out,
    output logic                    cp_ready,
    output logic                    cp_exception,
    
    // Debug Interface
    input  logic [ADDR_WIDTH-1:0]  debug_pc,
    input  logic [INST_WIDTH-1:0]  debug_instruction,
    input  logic [ADDR_WIDTH-1:0]  debug_mem_addr,
    input  logic [DATA_WIDTH-1:0]  debug_mem_data,
    input  logic                    debug_mem_write,
    input  logic                    debug_inst_valid,
    
    // Debug Control Outputs
    output logic                    debug_halt_request,
    output logic                    debug_single_step,
    output logic                    debug_breakpoint_hit,
    output logic                    debug_watchpoint_hit,
    
    // External Debug Interface
    input  logic                    external_debug_req,
    input  logic                    external_halt_req,
    output logic [DATA_WIDTH-1:0]  debug_status,
    output logic [ADDR_WIDTH-1:0]  debug_halt_pc
);

    // Debug register addresses
    typedef enum logic [11:0] {
        DBG_CTRL        = 12'h000,  // Debug control register
        DBG_STATUS      = 12'h001,  // Debug status register
        DBG_PC          = 12'h002,  // Current PC
        DBG_INST        = 12'h003,  // Current instruction
        DBG_BP_CTRL     = 12'h010,  // Breakpoint control
        DBG_BP_ADDR_BASE = 12'h020, // Breakpoint addresses start
        DBG_WP_CTRL     = 12'h030,  // Watchpoint control
        DBG_WP_ADDR_BASE = 12'h040, // Watchpoint addresses start
        DBG_WP_DATA_BASE = 12'h050, // Watchpoint data start
        DBG_PERF_CTR_BASE = 12'h100, // Performance counters start
        DBG_TRACE_CTRL  = 12'h200,  // Trace control
        DBG_TRACE_DATA  = 12'h201   // Trace data
    } dbg_reg_addr_t;
    
    // Instruction decode
    logic [6:0]  opcode;
    logic [2:0]  funct3;
    logic [11:0] csr_addr;
    logic [4:0]  rs1, rd;
    
    assign opcode = cp_instruction[6:0];
    assign funct3 = cp_instruction[14:12];
    assign csr_addr = cp_instruction[31:20];
    assign rs1 = cp_instruction[19:15];
    assign rd = cp_instruction[11:7];
    
    // Debug control registers
    logic [DATA_WIDTH-1:0] dbg_ctrl_reg;
    logic [DATA_WIDTH-1:0] dbg_status_reg;
    logic [DATA_WIDTH-1:0] dbg_pc_reg;
    logic [DATA_WIDTH-1:0] dbg_inst_reg;
    
    // Breakpoint registers
    logic [NUM_BREAKPOINTS-1:0] bp_enable;
    logic [ADDR_WIDTH-1:0] bp_addresses [NUM_BREAKPOINTS-1:0];
    logic [NUM_BREAKPOINTS-1:0] bp_hit;
    
    // Watchpoint registers
    logic [NUM_WATCHPOINTS-1:0] wp_enable;
    logic [NUM_WATCHPOINTS-1:0] wp_read_enable;
    logic [NUM_WATCHPOINTS-1:0] wp_write_enable;
    logic [ADDR_WIDTH-1:0] wp_addresses [NUM_WATCHPOINTS-1:0];
    logic [DATA_WIDTH-1:0] wp_data_values [NUM_WATCHPOINTS-1:0];
    logic [DATA_WIDTH-1:0] wp_data_masks [NUM_WATCHPOINTS-1:0];
    logic [NUM_WATCHPOINTS-1:0] wp_hit;
    
    // Performance counters
    logic [DATA_WIDTH-1:0] perf_cycle_count;
    logic [DATA_WIDTH-1:0] perf_inst_count;
    logic [DATA_WIDTH-1:0] perf_branch_count;
    logic [DATA_WIDTH-1:0] perf_cache_miss_count;
    
    // Trace buffer - using separate arrays instead of struct array for Icarus compatibility
    logic [ADDR_WIDTH-1:0]  trace_pc [TRACE_BUFFER_SIZE-1:0];
    logic [INST_WIDTH-1:0]  trace_instruction [TRACE_BUFFER_SIZE-1:0];
    logic [ADDR_WIDTH-1:0]  trace_mem_addr [TRACE_BUFFER_SIZE-1:0];
    logic [DATA_WIDTH-1:0]  trace_mem_data [TRACE_BUFFER_SIZE-1:0];
    logic                   trace_mem_write [TRACE_BUFFER_SIZE-1:0];
    logic [63:0]            trace_timestamp_buf [TRACE_BUFFER_SIZE-1:0];
    logic [$clog2(TRACE_BUFFER_SIZE)-1:0] trace_write_ptr;
    logic [$clog2(TRACE_BUFFER_SIZE)-1:0] trace_read_ptr;
    logic trace_enable;
    logic trace_full;
    logic trace_overflow;
    logic [63:0] trace_timestamp;
    
    // Debug state machine
    typedef enum logic [2:0] {
        DEBUG_RUNNING,
        DEBUG_HALTED,
        DEBUG_SINGLE_STEP,
        DEBUG_BREAKPOINT,
        DEBUG_WATCHPOINT
    } debug_state_t;
    
    debug_state_t debug_state;
    logic debug_halt_internal;
    logic debug_resume_req;
    logic debug_step_req;
    
    // Detect debug instructions
    logic is_debug_instruction;
    assign is_debug_instruction = cp_enable && (opcode == 7'b1110011) && (funct3 != 3'b000);
    
    // Breakpoint detection
    always_comb begin
        bp_hit = '0;
        for (int i = 0; i < NUM_BREAKPOINTS; i++) begin
            if (bp_enable[i] && (debug_pc == bp_addresses[i])) begin
                bp_hit[i] = 1'b1;
            end
        end
    end
    
    // Watchpoint detection
    always_comb begin
        wp_hit = '0;
        for (int i = 0; i < NUM_WATCHPOINTS; i++) begin
            if (wp_enable[i] && (debug_mem_addr == wp_addresses[i])) begin
                begin
                    logic data_match;
                    data_match = ((debug_mem_data & wp_data_masks[i]) == 
                                               (wp_data_values[i] & wp_data_masks[i]));
                    if ((wp_read_enable[i] && !debug_mem_write) ||
                        (wp_write_enable[i] && debug_mem_write)) begin
                        if (wp_data_masks[i] == '0 || data_match) begin
                            wp_hit[i] = 1'b1;
                        end
                    end
                end
            end
        end
    end
    
    // Debug state management
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            debug_state <= DEBUG_RUNNING;
            debug_halt_internal <= 1'b0;
        end else begin
            case (debug_state)
                DEBUG_RUNNING: begin
                    if (external_halt_req || (|bp_hit) || (|wp_hit)) begin
                        debug_state <= DEBUG_HALTED;
                        debug_halt_internal <= 1'b1;
                    end else if (debug_step_req) begin
                        debug_state <= DEBUG_SINGLE_STEP;
                    end
                end
                DEBUG_HALTED: begin
                    if (debug_resume_req) begin
                        debug_state <= DEBUG_RUNNING;
                        debug_halt_internal <= 1'b0;
                    end else if (debug_step_req) begin
                        debug_state <= DEBUG_SINGLE_STEP;
                    end
                end
                DEBUG_SINGLE_STEP: begin
                    // Execute one instruction then halt
                    debug_state <= DEBUG_HALTED;
                    debug_halt_internal <= 1'b1;
                end
                default: begin
                    debug_state <= DEBUG_RUNNING;
                end
            endcase
        end
    end
    
    // Performance counter updates
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            perf_cycle_count <= '0;
            perf_inst_count <= '0;
            perf_branch_count <= '0;
            perf_cache_miss_count <= '0;
        end else begin
            perf_cycle_count <= perf_cycle_count + 1;
            if (debug_inst_valid) begin
                perf_inst_count <= perf_inst_count + 1;
                // Count branches (simplified detection)
                if (debug_instruction[6:0] == 7'b1100011 || // Branch instructions
                    debug_instruction[6:0] == 7'b1101111 || // JAL
                    debug_instruction[6:0] == 7'b1100111) begin // JALR
                    perf_branch_count <= perf_branch_count + 1;
                end
            end
        end
    end
    
    // Trace buffer management
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            trace_write_ptr <= '0;
            trace_read_ptr <= '0;
            trace_enable <= 1'b0;
            trace_overflow <= 1'b0;
            trace_timestamp <= '0;
        end else begin
            trace_timestamp <= trace_timestamp + 1;
            
            if (trace_enable && debug_inst_valid) begin
                trace_pc[trace_write_ptr] <= debug_pc;
                trace_instruction[trace_write_ptr] <= debug_instruction;
                trace_mem_addr[trace_write_ptr] <= debug_mem_addr;
                trace_mem_data[trace_write_ptr] <= debug_mem_data;
                trace_mem_write[trace_write_ptr] <= debug_mem_write;
                trace_timestamp_buf[trace_write_ptr] <= trace_timestamp;
                
                if (trace_write_ptr == TRACE_BUFFER_SIZE - 1) begin
                    trace_write_ptr <= '0;
                    if (trace_read_ptr == 0) begin
                        trace_overflow <= 1'b1;
                    end
                end else begin
                    trace_write_ptr <= trace_write_ptr + 1;
                end
            end
        end
    end
    
    // Register read/write logic
    logic [DATA_WIDTH-1:0] reg_read_data;
    logic reg_write_enable;
    logic [DATA_WIDTH-1:0] reg_write_data;
    
    always_comb begin
        reg_read_data = '0;
        reg_write_enable = 1'b0;
        reg_write_data = cp_data_in;
        debug_resume_req = 1'b0;
        debug_step_req = 1'b0;
        
        if (is_debug_instruction) begin
            if (funct3 == 3'b001 || funct3 == 3'b010 || funct3 == 3'b011) begin // CSR operations
                case (csr_addr)
                    DBG_CTRL: begin
                        reg_read_data = dbg_ctrl_reg;
                        if (funct3 == 3'b001) begin // CSRRW
                            reg_write_enable = 1'b1;
                            debug_resume_req = reg_write_data[0];
                            debug_step_req = reg_write_data[1];
                        end
                    end
                    DBG_STATUS: begin
                        reg_read_data = dbg_status_reg;
                    end
                    DBG_PC: begin
                        reg_read_data = debug_pc;
                    end
                    DBG_TRACE_CTRL: begin
                        reg_read_data = {trace_overflow, trace_full, 62'b0} | trace_enable;
                        if (funct3 == 3'b001) begin
                            reg_write_enable = 1'b1;
                        end
                    end
                    DBG_TRACE_DATA: begin
                        if (trace_read_ptr != trace_write_ptr) begin
                            reg_read_data = trace_pc[trace_read_ptr];
                        end
                    end
                    default: begin
                        // Handle breakpoint and watchpoint registers
                        if (csr_addr >= DBG_BP_ADDR_BASE && csr_addr < DBG_BP_ADDR_BASE + NUM_BREAKPOINTS) begin
                            begin
                                logic [3:0] bp_idx;
                                bp_idx = csr_addr[3:0];
                                reg_read_data = bp_addresses[bp_idx];
                                if (funct3 == 3'b001) begin
                                    reg_write_enable = 1'b1;
                                end
                            end
                        end
                    end
                endcase
            end
        end
    end
    
    // Register updates
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            dbg_ctrl_reg <= '0;
            dbg_status_reg <= '0;
            trace_enable <= 1'b0;
            bp_enable <= '0;
            wp_enable <= '0;
            for (int i = 0; i < NUM_BREAKPOINTS; i++) begin
                bp_addresses[i] <= '0;
            end
            for (int i = 0; i < NUM_WATCHPOINTS; i++) begin
                wp_addresses[i] <= '0;
                wp_data_values[i] <= '0;
                wp_data_masks[i] <= '0;
            end
        end else begin
            // Update status register
            dbg_status_reg <= {
                58'b0,
                debug_state == DEBUG_HALTED,    // [5] Halted
                (|wp_hit),                      // [4] Watchpoint hit
                (|bp_hit),                      // [3] Breakpoint hit
                debug_state == DEBUG_SINGLE_STEP, // [2] Single step
                external_debug_req,             // [1] External debug request
                debug_state != DEBUG_RUNNING    // [0] Debug mode
            };
            
            if (reg_write_enable && is_debug_instruction) begin
                case (csr_addr)
                    DBG_CTRL: begin
                        dbg_ctrl_reg <= reg_write_data;
                    end
                    DBG_TRACE_CTRL: begin
                        trace_enable <= reg_write_data[0];
                    end
                    default: begin
                        if (csr_addr >= DBG_BP_ADDR_BASE && csr_addr < DBG_BP_ADDR_BASE + NUM_BREAKPOINTS) begin
                            begin
                                logic [3:0] bp_idx;
                                bp_idx = csr_addr[3:0];
                                bp_addresses[bp_idx] <= reg_write_data[ADDR_WIDTH-1:0];
                                bp_enable[bp_idx] <= 1'b1;
                            end
                        end
                    end
                endcase
            end
        end
    end
    
    // Output assignments
    assign cp_data_out = reg_read_data;
    assign cp_ready = 1'b1; // Debug operations complete immediately
    assign cp_exception = 1'b0; // No exceptions for debug operations
    
    assign debug_halt_request = debug_halt_internal;
    assign debug_single_step = (debug_state == DEBUG_SINGLE_STEP);
    assign debug_breakpoint_hit = (|bp_hit);
    assign debug_watchpoint_hit = (|wp_hit);
    assign debug_status = dbg_status_reg;
    assign debug_halt_pc = debug_pc;

endmodule

// Coprocessor FPU FSM
// Finite State Machine for Floating Point Unit operations

module coprocessor_fpu_fsm #(
    parameter DATA_WIDTH = 64
)(
    input  logic                    clk,
    input  logic                    rst_n,
    
    // Control Interface
    input  logic                    fpu_start,
    input  logic [4:0]              fpu_operation,
    input  logic [1:0]              fpu_format,
    output logic                    fpu_ready,
    output logic                    fpu_busy,
    output logic                    fpu_done,
    
    // Pipeline Control
    output logic                    stage_decode_en,
    output logic                    stage_unpack_en,
    output logic                    stage_execute_en,
    output logic                    stage_normalize_en,
    output logic                    stage_round_en,
    output logic                    stage_pack_en,
    
    // Exception Handling
    input  logic                    exception_detected,
    output logic                    exception_handled,
    
    // Cycle Counter
    output logic [4:0]              cycle_count,
    input  logic [4:0]              required_cycles
);

    // FSM States
    typedef enum logic [3:0] {
        FPU_IDLE        = 4'b0000,
        FPU_DECODE      = 4'b0001,
        FPU_UNPACK      = 4'b0010,
        FPU_EXECUTE     = 4'b0011,
        FPU_NORMALIZE   = 4'b0100,
        FPU_ROUND       = 4'b0101,
        FPU_PACK        = 4'b0110,
        FPU_COMPLETE    = 4'b0111,
        FPU_EXCEPTION   = 4'b1000,
        FPU_STALL       = 4'b1001
    } fpu_state_t;
    
    fpu_state_t current_state, next_state;
    
    // Internal counters and flags
    logic [4:0] cycle_counter;
    logic       operation_complete;
    logic       multi_cycle_op;
    
    // Determine if operation is multi-cycle
    always_comb begin
        multi_cycle_op = 1'b0;
        case (fpu_operation)
            5'b00011: multi_cycle_op = 1'b1; // DIV
            5'b00100: multi_cycle_op = 1'b1; // SQRT
            5'b00101,
            5'b00110,
            5'b00111,
            5'b01000: multi_cycle_op = 1'b1; // FMADD operations
            default:  multi_cycle_op = 1'b0;
        endcase
    end
    
    // State register
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            current_state <= FPU_IDLE;
            cycle_counter <= 5'b0;
        end else begin
            current_state <= next_state;
            
            if (current_state == FPU_EXECUTE) begin
                cycle_counter <= cycle_counter + 1;
            end else begin
                cycle_counter <= 5'b0;
            end
        end
    end
    
    // Next state logic
    always_comb begin
        next_state = current_state;
        operation_complete = (cycle_counter >= required_cycles);
        
        case (current_state)
            FPU_IDLE: begin
                if (fpu_start) begin
                    next_state = FPU_DECODE;
                end
            end
            
            FPU_DECODE: begin
                if (exception_detected) begin
                    next_state = FPU_EXCEPTION;
                end else begin
                    next_state = FPU_UNPACK;
                end
            end
            
            FPU_UNPACK: begin
                if (exception_detected) begin
                    next_state = FPU_EXCEPTION;
                end else begin
                    next_state = FPU_EXECUTE;
                end
            end
            
            FPU_EXECUTE: begin
                if (exception_detected) begin
                    next_state = FPU_EXCEPTION;
                end else if (multi_cycle_op && !operation_complete) begin
                    next_state = FPU_EXECUTE; // Stay in execute
                end else begin
                    next_state = FPU_NORMALIZE;
                end
            end
            
            FPU_NORMALIZE: begin
                if (exception_detected) begin
                    next_state = FPU_EXCEPTION;
                end else begin
                    next_state = FPU_ROUND;
                end
            end
            
            FPU_ROUND: begin
                if (exception_detected) begin
                    next_state = FPU_EXCEPTION;
                end else begin
                    next_state = FPU_PACK;
                end
            end
            
            FPU_PACK: begin
                next_state = FPU_COMPLETE;
            end
            
            FPU_COMPLETE: begin
                next_state = FPU_IDLE;
            end
            
            FPU_EXCEPTION: begin
                next_state = FPU_IDLE;
            end
            
            FPU_STALL: begin
                // Future use for pipeline stalls
                next_state = FPU_IDLE;
            end
            
            default: begin
                next_state = FPU_IDLE;
            end
        endcase
    end
    
    // Output control signals
    always_comb begin
        // Default values
        stage_decode_en = 1'b0;
        stage_unpack_en = 1'b0;
        stage_execute_en = 1'b0;
        stage_normalize_en = 1'b0;
        stage_round_en = 1'b0;
        stage_pack_en = 1'b0;
        fpu_ready = 1'b0;
        fpu_busy = 1'b0;
        fpu_done = 1'b0;
        exception_handled = 1'b0;
        
        case (current_state)
            FPU_IDLE: begin
                fpu_ready = 1'b1;
            end
            
            FPU_DECODE: begin
                stage_decode_en = 1'b1;
                fpu_busy = 1'b1;
            end
            
            FPU_UNPACK: begin
                stage_unpack_en = 1'b1;
                fpu_busy = 1'b1;
            end
            
            FPU_EXECUTE: begin
                stage_execute_en = 1'b1;
                fpu_busy = 1'b1;
            end
            
            FPU_NORMALIZE: begin
                stage_normalize_en = 1'b1;
                fpu_busy = 1'b1;
            end
            
            FPU_ROUND: begin
                stage_round_en = 1'b1;
                fpu_busy = 1'b1;
            end
            
            FPU_PACK: begin
                stage_pack_en = 1'b1;
                fpu_busy = 1'b1;
            end
            
            FPU_COMPLETE: begin
                fpu_done = 1'b1;
            end
            
            FPU_EXCEPTION: begin
                exception_handled = 1'b1;
            end
            
            default: begin
                fpu_ready = 1'b1;
            end
        endcase
    end
    
    // Cycle count output
    assign cycle_count = cycle_counter;

endmodule

// Coprocessor FPU
// Floating Point Unit for coprocessor operations

module coprocessor_fpu #(
    parameter DATA_WIDTH = 64,
    parameter ADDR_WIDTH = 64,
    parameter INST_WIDTH = 32
)(
    input  logic                    clk,
    input  logic                    rst_n,
    
    // Coprocessor Interface
    input  logic                    cp_enable,
    input  logic [INST_WIDTH-1:0]  cp_instruction,
    input  logic [DATA_WIDTH-1:0]  cp_data_in,
    output logic [DATA_WIDTH-1:0]  cp_data_out,
    output logic                    cp_ready,
    output logic                    cp_exception,
    
    // FPU Register File Interface
    output logic                    fp_reg_write,
    output logic [4:0]              fp_reg_waddr,
    output logic [DATA_WIDTH-1:0]   fp_reg_wdata,
    output logic [4:0]              fp_reg_raddr1,
    output logic [4:0]              fp_reg_raddr2,
    output logic [4:0]              fp_reg_raddr3,
    input  logic [DATA_WIDTH-1:0]   fp_reg_rdata1,
    input  logic [DATA_WIDTH-1:0]   fp_reg_rdata2,
    input  logic [DATA_WIDTH-1:0]   fp_reg_rdata3,
    
    // Status and Control
    output logic [4:0]              fpu_flags,
    output logic                    fpu_busy
);

    // Instruction decode
    logic [6:0]  opcode;
    logic [4:0]  rd, rs1, rs2, rs3;
    logic [2:0]  funct3;
    logic [6:0]  funct7;
    logic [1:0]  fmt;
    logic [2:0]  rm;
    
    assign opcode = cp_instruction[6:0];
    assign rd = cp_instruction[11:7];
    assign funct3 = cp_instruction[14:12];
    assign rs1 = cp_instruction[19:15];
    assign rs2 = cp_instruction[24:20];
    assign funct7 = cp_instruction[31:25];
    assign rs3 = cp_instruction[31:27];
    assign fmt = cp_instruction[26:25];
    assign rm = cp_instruction[14:12];
    
    // FPU operation encoding
    logic [4:0] fpu_operation;
    logic [1:0] fpu_format;
    logic [2:0] fpu_rounding;
    logic       fpu_start;
    logic       fpu_done;
    logic       fpu_ready_internal;
    logic       exception_detected;
    
    // FSM interface
    logic       stage_decode_en;
    logic       stage_unpack_en;
    logic       stage_execute_en;
    logic       stage_normalize_en;
    logic       stage_round_en;
    logic       stage_pack_en;
    logic [4:0] cycle_count;
    logic [4:0] required_cycles;
    
    // Operands and results
    logic [DATA_WIDTH-1:0] operand_a, operand_b, operand_c;
    logic [DATA_WIDTH-1:0] fpu_result;
    logic                  result_valid;
    
    // Exception flags
    logic flag_invalid, flag_div_zero, flag_overflow, flag_underflow, flag_inexact;
    
    // Instruction decoding
    always_comb begin
        fpu_operation = 5'b0;
        fpu_format = fmt;
        fpu_rounding = rm;
        fpu_start = 1'b0;
        
        if (cp_enable) begin
            case (opcode)
                7'b1010011: begin // FP_OP
                    fpu_start = 1'b1;
                    case (funct7)
                        7'b0000000: fpu_operation = 5'b00000; // FADD
                        7'b0000100: fpu_operation = 5'b00001; // FSUB
                        7'b0001000: fpu_operation = 5'b00010; // FMUL
                        7'b0001100: fpu_operation = 5'b00011; // FDIV
                        7'b0101100: fpu_operation = 5'b00100; // FSQRT
                        7'b0010000: begin // FSGNJ
                            case (funct3)
                                3'b000: fpu_operation = 5'b01011; // FSGNJ
                                3'b001: fpu_operation = 5'b01100; // FSGNJN
                                3'b010: fpu_operation = 5'b01101; // FSGNJX
                            endcase
                        end
                        7'b0010100: begin // FMIN/FMAX
                            case (funct3)
                                3'b000: fpu_operation = 5'b01001; // FMIN
                                3'b001: fpu_operation = 5'b01010; // FMAX
                            endcase
                        end
                        7'b1010000: begin // FP Compare
                            case (funct3)
                                3'b010: fpu_operation = 5'b01110; // FEQ
                                3'b001: fpu_operation = 5'b01111; // FLT
                                3'b000: fpu_operation = 5'b10000; // FLE
                            endcase
                        end
                        7'b1100000: begin // FP to INT
                            case (rs2)
                                5'b00000: fpu_operation = 5'b10001; // FCVT.W.S/D
                                5'b00001: fpu_operation = 5'b10010; // FCVT.WU.S/D
                                5'b00010: fpu_operation = 5'b10011; // FCVT.L.S/D
                                5'b00011: fpu_operation = 5'b10100; // FCVT.LU.S/D
                            endcase
                        end
                        7'b1101000: begin // INT to FP (single)
                            case (rs2)
                                5'b00000: fpu_operation = 5'b10101; // FCVT.S.W
                                5'b00001: fpu_operation = 5'b10101; // FCVT.S.WU
                                5'b00010: fpu_operation = 5'b10101; // FCVT.S.L
                                5'b00011: fpu_operation = 5'b10101; // FCVT.S.LU
                            endcase
                        end
                        7'b1101001: begin // INT to FP (double)
                            case (rs2)
                                5'b00000: fpu_operation = 5'b10110; // FCVT.D.W
                                5'b00001: fpu_operation = 5'b10110; // FCVT.D.WU
                                5'b00010: fpu_operation = 5'b10110; // FCVT.D.L
                                5'b00011: fpu_operation = 5'b10110; // FCVT.D.LU
                            endcase
                        end
                        7'b0100000: begin // FP conversion
                            if (rs2 == 5'b00001) begin
                                fpu_operation = 5'b10111; // FCVT.S.D
                            end
                        end
                        7'b0100001: begin // FP conversion
                            if (rs2 == 5'b00000) begin
                                fpu_operation = 5'b11000; // FCVT.D.S
                            end
                        end
                        7'b1110000: fpu_operation = 5'b11001; // FCLASS
                        7'b1111000: fpu_operation = 5'b11010; // FMV
                        default: fpu_operation = 5'b0;
                    endcase
                end
                7'b1000011: begin // FMADD
                    fpu_start = 1'b1;
                    fpu_operation = 5'b00101;
                end
                7'b1000111: begin // FMSUB
                    fpu_start = 1'b1;
                    fpu_operation = 5'b00110;
                end
                7'b1001011: begin // FNMSUB
                    fpu_start = 1'b1;
                    fpu_operation = 5'b00111;
                end
                7'b1001111: begin // FNMADD
                    fpu_start = 1'b1;
                    fpu_operation = 5'b01000;
                end
                default: begin
                    fpu_start = 1'b0;
                end
            endcase
        end
    end
    
    // Determine required cycles for operation
    always_comb begin
        case (fpu_operation)
            5'b00000, 5'b00001: required_cycles = 5'd3;  // ADD/SUB
            5'b00010:           required_cycles = 5'd4;  // MUL
            5'b00011:           required_cycles = 5'd16; // DIV
            5'b00100:           required_cycles = 5'd20; // SQRT
            5'b00101, 5'b00110,
            5'b00111, 5'b01000: required_cycles = 5'd5;  // FMADD operations
            5'b10001, 5'b10010,
            5'b10011, 5'b10100,
            5'b10101, 5'b10110,
            5'b10111, 5'b11000: required_cycles = 5'd2;  // Conversions
            default:            required_cycles = 5'd1;  // Single cycle ops
        endcase
    end
    
    // Operand selection
    always_comb begin
        operand_a = fp_reg_rdata1;
        operand_b = fp_reg_rdata2;
        operand_c = fp_reg_rdata3;
        
        // For load/store operations, use CPU data
        if (opcode == 7'b0000111 || opcode == 7'b0100111) begin
            operand_a = cp_data_in;
        end
        
        // For move operations from integer
        if (funct7 == 7'b1111000 && rs2[0]) begin
            operand_a = cp_data_in;
        end
    end
    
    // FPU FSM instantiation
    coprocessor_fpu_fsm fpu_fsm (
        .clk(clk),
        .rst_n(rst_n),
        .fpu_start(fpu_start),
        .fpu_operation(fpu_operation),
        .fpu_format(fpu_format),
        .fpu_ready(fpu_ready_internal),
        .fpu_busy(fpu_busy),
        .fpu_done(fpu_done),
        .stage_decode_en(stage_decode_en),
        .stage_unpack_en(stage_unpack_en),
        .stage_execute_en(stage_execute_en),
        .stage_normalize_en(stage_normalize_en),
        .stage_round_en(stage_round_en),
        .stage_pack_en(stage_pack_en),
        .exception_detected(exception_detected),
        .exception_handled(),
        .cycle_count(cycle_count),
        .required_cycles(required_cycles)
    );
    
    // Simplified FPU execution core
    logic [DATA_WIDTH-1:0] exec_result;
    logic exec_valid;
    
    always_comb begin
        exec_result = operand_a; // Default passthrough
        exec_valid = stage_pack_en;
        exception_detected = 1'b0;
        
        // Simplified operation execution
        if (stage_execute_en) begin
            case (fpu_operation)
                5'b00000: begin // FADD
                    // Simplified: would need proper IEEE 754 addition
                    exec_result = operand_a;
                end
                5'b00001: begin // FSUB
                    exec_result = operand_a;
                end
                5'b00010: begin // FMUL
                    exec_result = operand_a;
                end
                5'b00011: begin // FDIV
                    exec_result = operand_a;
                    if (operand_b == 64'b0) begin
                        exception_detected = 1'b1;
                    end
                end
                5'b01110: begin // FEQ
                    exec_result = (operand_a == operand_b) ? 64'b1 : 64'b0;
                end
                5'b01111: begin // FLT
                    exec_result = (operand_a < operand_b) ? 64'b1 : 64'b0;
                end
                5'b10000: begin // FLE
                    exec_result = (operand_a <= operand_b) ? 64'b1 : 64'b0;
                end
                5'b11010: begin // FMV
                    exec_result = operand_a;
                end
                default: begin
                    exec_result = operand_a;
                end
            endcase
        end
    end
    
    // Result capture
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            fpu_result <= 64'b0;
            result_valid <= 1'b0;
        end else begin
            if (exec_valid) begin
                fpu_result <= exec_result;
                result_valid <= 1'b1;
            end else if (fpu_done) begin
                result_valid <= 1'b0;
            end
        end
    end
    
    // Exception flag generation (simplified)
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            flag_invalid <= 1'b0;
            flag_div_zero <= 1'b0;
            flag_overflow <= 1'b0;
            flag_underflow <= 1'b0;
            flag_inexact <= 1'b0;
        end else begin
            if (exception_detected) begin
                flag_div_zero <= (fpu_operation == 5'b00011); // DIV
                flag_invalid <= 1'b1;
            end else if (fpu_done) begin
                flag_invalid <= 1'b0;
                flag_div_zero <= 1'b0;
                flag_overflow <= 1'b0;
                flag_underflow <= 1'b0;
                flag_inexact <= 1'b0;
            end
        end
    end
    
    // Register file connections
    assign fp_reg_raddr1 = rs1;
    assign fp_reg_raddr2 = rs2;
    assign fp_reg_raddr3 = rs3;
    assign fp_reg_write = fpu_done && (rd != 5'b0) && (opcode != 7'b0100111); // Not store
    assign fp_reg_waddr = rd;
    assign fp_reg_wdata = fpu_result;
    
    // Output assignments
    assign cp_data_out = fpu_result;
    assign cp_ready = fpu_ready_internal;
    assign cp_exception = exception_detected;
    assign fpu_flags = {flag_invalid, flag_div_zero, flag_overflow, flag_underflow, flag_inexact};

endmodule

// Coprocessor FSM
// Generic Finite State Machine for coprocessor operations

module coprocessor_fsm #(
    parameter DATA_WIDTH = 64,
    parameter STATE_WIDTH = 4,
    parameter OP_WIDTH = 5
)(
    input  logic                    clk,
    input  logic                    rst_n,
    
    // Control Interface
    input  logic                    cp_start,
    input  logic [OP_WIDTH-1:0]     cp_operation,
    input  logic                    cp_stall,
    output logic                    cp_ready,
    output logic                    cp_busy,
    output logic                    cp_done,
    
    // Pipeline Stage Control
    output logic                    stage_fetch_en,
    output logic                    stage_decode_en,
    output logic                    stage_execute_en,
    output logic                    stage_writeback_en,
    
    // Exception Handling
    input  logic                    exception_request,
    input  logic [3:0]              exception_code,
    output logic                    exception_active,
    output logic                    exception_handled,
    
    // Multi-cycle Operation Support
    input  logic [7:0]              required_cycles,
    output logic [7:0]              current_cycle,
    output logic                    operation_complete,
    
    // Debug Interface
    output logic [STATE_WIDTH-1:0] current_state_debug,
    output logic [STATE_WIDTH-1:0] next_state_debug
);

    // FSM States
    typedef enum logic [STATE_WIDTH-1:0] {
        CP_IDLE         = 4'b0000,
        CP_FETCH        = 4'b0001,
        CP_DECODE       = 4'b0010,
        CP_EXECUTE      = 4'b0011,
        CP_WRITEBACK    = 4'b0100,
        CP_COMPLETE     = 4'b0101,
        CP_EXCEPTION    = 4'b0110,
        CP_STALL        = 4'b0111,
        CP_FLUSH        = 4'b1000,
        CP_RESET        = 4'b1001
    } cp_state_t;
    
    cp_state_t current_state, next_state;
    
    // Internal registers
    logic [7:0]  cycle_counter;
    logic [OP_WIDTH-1:0] operation_reg;
    logic        multi_cycle_operation;
    logic        exception_pending;
    logic [3:0]  exception_code_reg;
    
    // Operation classification
    always_comb begin
        multi_cycle_operation = 1'b0;
        case (cp_operation)
            5'b00011,  // Division
            5'b00100,  // Square root
            5'b00101,  // Multiply-add
            5'b00110,  // Multiply-sub
            5'b00111,  // Negative multiply-add
            5'b01000,  // Negative multiply-sub
            5'b10000,  // Load/Store operations
            5'b10001,  // Memory operations
            5'b11000,  // System operations
            5'b11001:  // Debug operations
                multi_cycle_operation = 1'b1;
            default:
                multi_cycle_operation = 1'b0;
        endcase
    end
    
    // State register
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            current_state <= CP_IDLE;
            cycle_counter <= 8'b0;
            operation_reg <= '0;
            exception_pending <= 1'b0;
            exception_code_reg <= 4'b0;
        end else begin
            current_state <= next_state;
            
            // Cycle counter management
            if (current_state == CP_EXECUTE) begin
                cycle_counter <= cycle_counter + 1;
            end else begin
                cycle_counter <= 8'b0;
            end
            
            // Operation register
            if (current_state == CP_DECODE) begin
                operation_reg <= cp_operation;
            end
            
            // Exception handling
            if (exception_request && current_state != CP_EXCEPTION) begin
                exception_pending <= 1'b1;
                exception_code_reg <= exception_code;
            end else if (current_state == CP_EXCEPTION) begin
                exception_pending <= 1'b0;
            end
        end
    end
    
    // Next state logic
    always_comb begin
        next_state = current_state;
        operation_complete = (cycle_counter >= required_cycles);
        
        case (current_state)
            CP_IDLE: begin
                if (exception_request || exception_pending) begin
                    next_state = CP_EXCEPTION;
                end else if (cp_start) begin
                    next_state = CP_FETCH;
                end
            end
            
            CP_FETCH: begin
                if (exception_request || exception_pending) begin
                    next_state = CP_EXCEPTION;
                end else if (cp_stall) begin
                    next_state = CP_STALL;
                end else begin
                    next_state = CP_DECODE;
                end
            end
            
            CP_DECODE: begin
                if (exception_request || exception_pending) begin
                    next_state = CP_EXCEPTION;
                end else if (cp_stall) begin
                    next_state = CP_STALL;
                end else begin
                    next_state = CP_EXECUTE;
                end
            end
            
            CP_EXECUTE: begin
                if (exception_request || exception_pending) begin
                    next_state = CP_EXCEPTION;
                end else if (cp_stall) begin
                    next_state = CP_STALL;
                end else if (multi_cycle_operation && !operation_complete) begin
                    next_state = CP_EXECUTE; // Stay in execute
                end else begin
                    next_state = CP_WRITEBACK;
                end
            end
            
            CP_WRITEBACK: begin
                if (exception_request || exception_pending) begin
                    next_state = CP_EXCEPTION;
                end else if (cp_stall) begin
                    next_state = CP_STALL;
                end else begin
                    next_state = CP_COMPLETE;
                end
            end
            
            CP_COMPLETE: begin
                next_state = CP_IDLE;
            end
            
            CP_EXCEPTION: begin
                // Stay in exception state for one cycle
                next_state = CP_IDLE;
            end
            
            CP_STALL: begin
                if (exception_request || exception_pending) begin
                    next_state = CP_EXCEPTION;
                end else if (!cp_stall) begin
                    // Return to previous state logic
                    case (operation_reg)
                        default: next_state = CP_EXECUTE;
                    endcase
                end
            end
            
            CP_FLUSH: begin
                next_state = CP_IDLE;
            end
            
            CP_RESET: begin
                next_state = CP_IDLE;
            end
            
            default: begin
                next_state = CP_IDLE;
            end
        endcase
    end
    
    // Output control signals
    always_comb begin
        // Default values
        stage_fetch_en = 1'b0;
        stage_decode_en = 1'b0;
        stage_execute_en = 1'b0;
        stage_writeback_en = 1'b0;
        cp_ready = 1'b0;
        cp_busy = 1'b0;
        cp_done = 1'b0;
        exception_active = 1'b0;
        exception_handled = 1'b0;
        
        case (current_state)
            CP_IDLE: begin
                cp_ready = 1'b1;
            end
            
            CP_FETCH: begin
                stage_fetch_en = 1'b1;
                cp_busy = 1'b1;
            end
            
            CP_DECODE: begin
                stage_decode_en = 1'b1;
                cp_busy = 1'b1;
            end
            
            CP_EXECUTE: begin
                stage_execute_en = 1'b1;
                cp_busy = 1'b1;
            end
            
            CP_WRITEBACK: begin
                stage_writeback_en = 1'b1;
                cp_busy = 1'b1;
            end
            
            CP_COMPLETE: begin
                cp_done = 1'b1;
            end
            
            CP_EXCEPTION: begin
                exception_active = 1'b1;
                exception_handled = 1'b1;
            end
            
            CP_STALL: begin
                cp_busy = 1'b1;
            end
            
            CP_FLUSH: begin
                // Flush state - no enables
            end
            
            CP_RESET: begin
                // Reset state - no enables
            end
            
            default: begin
                cp_ready = 1'b1;
            end
        endcase
    end
    
    // Cycle counter output
    assign current_cycle = cycle_counter;
    
    // Debug outputs
    assign current_state_debug = current_state;
    assign next_state_debug = next_state;

endmodule

// Coprocessor Integer ALU
// Specialized ALU for coprocessor integer operations

module coprocessor_int_alu #(
    parameter DATA_WIDTH = 64,
    parameter ADDR_WIDTH = 64
)(
    input  logic                    clk,
    input  logic                    rst_n,
    
    // Control Interface
    input  logic                    alu_enable,
    input  logic [4:0]              alu_operation,
    input  logic [2:0]              alu_format,
    
    // Data Interface
    input  logic [DATA_WIDTH-1:0]  operand_a,
    input  logic [DATA_WIDTH-1:0]  operand_b,
    input  logic [DATA_WIDTH-1:0]  operand_c,
    output logic [DATA_WIDTH-1:0]  result,
    output logic                    result_valid,
    
    // Status Flags
    output logic                    zero_flag,
    output logic                    negative_flag,
    output logic                    carry_flag,
    output logic                    overflow_flag,
    output logic                    parity_flag,
    
    // Control Outputs
    output logic                    alu_ready,
    output logic                    alu_busy
);

    // ALU Operation Codes
    typedef enum logic [4:0] {
        ALU_ADD     = 5'b00000,
        ALU_SUB     = 5'b00001,
        ALU_AND     = 5'b00010,
        ALU_OR      = 5'b00011,
        ALU_XOR     = 5'b00100,
        ALU_SLL     = 5'b00101,  // Shift left logical
        ALU_SRL     = 5'b00110,  // Shift right logical
        ALU_SRA     = 5'b00111,  // Shift right arithmetic
        ALU_SLT     = 5'b01000,  // Set less than
        ALU_SLTU    = 5'b01001,  // Set less than unsigned
        ALU_MUL     = 5'b01010,  // Multiply
        ALU_MULH    = 5'b01011,  // Multiply high
        ALU_MULHU   = 5'b01100,  // Multiply high unsigned
        ALU_MULHSU  = 5'b01101,  // Multiply high signed-unsigned
        ALU_DIV     = 5'b01110,  // Divide
        ALU_DIVU    = 5'b01111,  // Divide unsigned
        ALU_REM     = 5'b10000,  // Remainder
        ALU_REMU    = 5'b10001,  // Remainder unsigned
        ALU_MAX     = 5'b10010,  // Maximum
        ALU_MIN     = 5'b10011,  // Minimum
        ALU_MAXU    = 5'b10100,  // Maximum unsigned
        ALU_MINU    = 5'b10101,  // Minimum unsigned
        ALU_CLZ     = 5'b10110,  // Count leading zeros
        ALU_CTZ     = 5'b10111,  // Count trailing zeros
        ALU_PCNT    = 5'b11000,  // Population count
        ALU_BSWAP   = 5'b11001,  // Byte swap
        ALU_SEXT_B  = 5'b11010,  // Sign extend byte
        ALU_SEXT_H  = 5'b11011,  // Sign extend halfword
        ALU_ZEXT_B  = 5'b11100,  // Zero extend byte
        ALU_ZEXT_H  = 5'b11101,  // Zero extend halfword
        ALU_ROL     = 5'b11110,  // Rotate left
        ALU_ROR     = 5'b11111   // Rotate right
    } alu_op_t;
    
    // Format types
    typedef enum logic [2:0] {
        FMT_WORD    = 3'b000,    // 32-bit operation
        FMT_DWORD   = 3'b001,    // 64-bit operation
        FMT_BYTE    = 3'b010,    // 8-bit operation
        FMT_HWORD   = 3'b011,    // 16-bit operation
        FMT_SIGNED  = 3'b100,    // Signed operation
        FMT_UNSIGNED = 3'b101    // Unsigned operation
    } alu_fmt_t;
    
    // Internal signals
    logic [DATA_WIDTH-1:0]   alu_result;
    logic [DATA_WIDTH*2-1:0] extended_result;  // For multiply operations
    logic [5:0]              shift_amount;
    logic                    operation_done;
    logic                    multi_cycle_op;
    logic [3:0]              cycle_counter;
    
    // Status flag computation
    logic result_zero, result_negative, result_carry, result_overflow, result_parity;
    
    // Determine if operation is multi-cycle
    always_comb begin
        multi_cycle_op = 1'b0;
        case (alu_operation)
            ALU_MUL, ALU_MULH, ALU_MULHU, ALU_MULHSU,
            ALU_DIV, ALU_DIVU, ALU_REM, ALU_REMU:
                multi_cycle_op = 1'b1;
            default:
                multi_cycle_op = 1'b0;
        endcase
    end
    
    // Shift amount extraction
    always_comb begin
        if (alu_format == FMT_WORD) begin
            shift_amount = operand_b[4:0];  // 32-bit shifts use 5 bits
        end else begin
            shift_amount = operand_b[5:0];  // 64-bit shifts use 6 bits
        end
    end
    
    // Multi-cycle operation counter
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            cycle_counter <= 4'b0;
            operation_done <= 1'b0;
        end else begin
            if (alu_enable && multi_cycle_op) begin
                if (cycle_counter < 4'd8) begin // Max 8 cycles for complex ops
                    cycle_counter <= cycle_counter + 1;
                    operation_done <= 1'b0;
                end else begin
                    operation_done <= 1'b1;
                    cycle_counter <= 4'b0;
                end
            end else if (alu_enable) begin
                operation_done <= 1'b1;
                cycle_counter <= 4'b0;
            end else begin
                operation_done <= 1'b0;
                cycle_counter <= 4'b0;
            end
        end
    end
    
    // Main ALU logic
    always_comb begin
        alu_result = 64'b0;
        extended_result = 128'b0;
        result_carry = 1'b0;
        result_overflow = 1'b0;
        
        case (alu_operation)
            ALU_ADD: begin
                {result_carry, alu_result} = operand_a + operand_b;
                result_overflow = (operand_a[DATA_WIDTH-1] == operand_b[DATA_WIDTH-1]) &&
                                 (alu_result[DATA_WIDTH-1] != operand_a[DATA_WIDTH-1]);
            end
            
            ALU_SUB: begin
                {result_carry, alu_result} = operand_a - operand_b;
                result_overflow = (operand_a[DATA_WIDTH-1] != operand_b[DATA_WIDTH-1]) &&
                                 (alu_result[DATA_WIDTH-1] != operand_a[DATA_WIDTH-1]);
            end
            
            ALU_AND: begin
                alu_result = operand_a & operand_b;
            end
            
            ALU_OR: begin
                alu_result = operand_a | operand_b;
            end
            
            ALU_XOR: begin
                alu_result = operand_a ^ operand_b;
            end
            
            ALU_SLL: begin
                if (alu_format == FMT_WORD) begin
                    alu_result = {{32{1'b0}}, operand_a[31:0] << shift_amount[4:0]};
                end else begin
                    alu_result = operand_a << shift_amount;
                end
            end
            
            ALU_SRL: begin
                if (alu_format == FMT_WORD) begin
                    alu_result = {{32{1'b0}}, operand_a[31:0] >> shift_amount[4:0]};
                end else begin
                    alu_result = operand_a >> shift_amount;
                end
            end
            
            ALU_SRA: begin
                if (alu_format == FMT_WORD) begin
                    alu_result = {{32{operand_a[31]}}, $signed(operand_a[31:0]) >>> shift_amount[4:0]};
                end else begin
                    alu_result = $signed(operand_a) >>> shift_amount;
                end
            end
            
            ALU_SLT: begin
                alu_result = ($signed(operand_a) < $signed(operand_b)) ? 64'b1 : 64'b0;
            end
            
            ALU_SLTU: begin
                alu_result = (operand_a < operand_b) ? 64'b1 : 64'b0;
            end
            
            ALU_MUL: begin
                if (alu_format == FMT_WORD) begin
                    extended_result = $signed(operand_a[31:0]) * $signed(operand_b[31:0]);
                    alu_result = {{32{extended_result[31]}}, extended_result[31:0]};
                end else begin
                    extended_result = $signed(operand_a) * $signed(operand_b);
                    alu_result = extended_result[63:0];
                end
            end
            
            ALU_MULH: begin
                extended_result = $signed(operand_a) * $signed(operand_b);
                alu_result = extended_result[127:64];
            end
            
            ALU_MULHU: begin
                extended_result = operand_a * operand_b;
                alu_result = extended_result[127:64];
            end
            
            ALU_MULHSU: begin
                extended_result = $signed(operand_a) * operand_b;
                alu_result = extended_result[127:64];
            end
            
            ALU_DIV: begin
                if (operand_b != 64'b0) begin
                    alu_result = $signed(operand_a) / $signed(operand_b);
                end else begin
                    alu_result = 64'hFFFFFFFFFFFFFFFF; // Division by zero
                end
            end
            
            ALU_DIVU: begin
                if (operand_b != 64'b0) begin
                    alu_result = operand_a / operand_b;
                end else begin
                    alu_result = 64'hFFFFFFFFFFFFFFFF; // Division by zero
                end
            end
            
            ALU_REM: begin
                if (operand_b != 64'b0) begin
                    alu_result = $signed(operand_a) % $signed(operand_b);
                end else begin
                    alu_result = operand_a; // Remainder by zero
                end
            end
            
            ALU_REMU: begin
                if (operand_b != 64'b0) begin
                    alu_result = operand_a % operand_b;
                end else begin
                    alu_result = operand_a; // Remainder by zero
                end
            end
            
            ALU_MAX: begin
                alu_result = ($signed(operand_a) > $signed(operand_b)) ? operand_a : operand_b;
            end
            
            ALU_MIN: begin
                alu_result = ($signed(operand_a) < $signed(operand_b)) ? operand_a : operand_b;
            end
            
            ALU_MAXU: begin
                alu_result = (operand_a > operand_b) ? operand_a : operand_b;
            end
            
            ALU_MINU: begin
                alu_result = (operand_a < operand_b) ? operand_a : operand_b;
            end
            
            ALU_CLZ: begin // Count leading zeros
                alu_result = 64'b0;
                for (int i = 63; i >= 0; i--) begin
                    if (operand_a[i] == 1'b0) begin
                        alu_result = alu_result + 1;
                    end else begin
                        i = -1; // Exit loop
                    end
                end
            end
            
            ALU_CTZ: begin // Count trailing zeros
                alu_result = 64'b0;
                for (int i = 0; i < 64; i++) begin
                    if (operand_a[i] == 1'b0) begin
                        alu_result = alu_result + 1;
                    end else begin
                        i = 64; // Exit loop
                    end
                end
            end
            
            ALU_PCNT: begin // Population count
                alu_result = 64'b0;
                for (int i = 0; i < 64; i++) begin
                    alu_result = alu_result + operand_a[i];
                end
            end
            
            ALU_BSWAP: begin // Byte swap
                alu_result = {operand_a[7:0], operand_a[15:8], operand_a[23:16], operand_a[31:24],
                             operand_a[39:32], operand_a[47:40], operand_a[55:48], operand_a[63:56]};
            end
            
            ALU_SEXT_B: begin // Sign extend byte
                alu_result = {{56{operand_a[7]}}, operand_a[7:0]};
            end
            
            ALU_SEXT_H: begin // Sign extend halfword
                alu_result = {{48{operand_a[15]}}, operand_a[15:0]};
            end
            
            ALU_ZEXT_B: begin // Zero extend byte
                alu_result = {56'b0, operand_a[7:0]};
            end
            
            ALU_ZEXT_H: begin // Zero extend halfword
                alu_result = {48'b0, operand_a[15:0]};
            end
            
            ALU_ROL: begin // Rotate left
                alu_result = (operand_a << shift_amount) | (operand_a >> (64 - shift_amount));
            end
            
            ALU_ROR: begin // Rotate right
                alu_result = (operand_a >> shift_amount) | (operand_a << (64 - shift_amount));
            end
            
            default: begin
                alu_result = operand_a;
            end
        endcase
    end
    
    // Status flag computation
    always_comb begin
        result_zero = (alu_result == 64'b0);
        result_negative = alu_result[DATA_WIDTH-1];
        
        // Parity calculation (even parity)
        result_parity = 1'b0;
        for (int i = 0; i < 8; i++) begin
            result_parity = result_parity ^ alu_result[i];
        end
    end
    
    // Output assignments
    assign result = alu_result;
    assign result_valid = operation_done;
    assign alu_ready = !alu_enable || operation_done;
    assign alu_busy = alu_enable && !operation_done;
    
    // Status flags
    assign zero_flag = result_zero;
    assign negative_flag = result_negative;
    assign carry_flag = result_carry;
    assign overflow_flag = result_overflow;
    assign parity_flag = result_parity;

endmodule

// Coprocessor Interface
// Defines the interface between CPU and coprocessors for system operations

module coprocessor_interface #(
    parameter ADDR_WIDTH = 64,
    parameter DATA_WIDTH = 64,
    parameter INST_WIDTH = 32,
    parameter CP_NUM = 4  // Number of coprocessors
)(
    input  logic                    clk,
    input  logic                    rst_n,
    
    // CPU Interface
    input  logic                    cp_valid,        // Coprocessor instruction valid
    input  logic [INST_WIDTH-1:0]  cp_instruction,  // Coprocessor instruction
    input  logic [DATA_WIDTH-1:0]  cp_data_in,      // Data from CPU
    output logic [DATA_WIDTH-1:0]  cp_data_out,     // Data to CPU
    output logic                    cp_ready,        // Coprocessor ready
    output logic                    cp_exception,    // Exception occurred
    
    // Coprocessor Select
    input  logic [1:0]              cp_select,       // Which coprocessor (0-3)
    
    // Individual Coprocessor Interfaces
    output logic [CP_NUM-1:0]       cp_enable,       // Enable signals for each CP
    output logic [INST_WIDTH-1:0]   cp_inst_out,     // Instruction to selected CP
    output logic [DATA_WIDTH-1:0]   cp_data_to_cp,   // Data to selected CP
    input  logic [DATA_WIDTH-1:0]   cp_data_from_cp [CP_NUM-1:0], // Data from CPs
    input  logic [CP_NUM-1:0]       cp_ready_in,     // Ready signals from CPs
    input  logic [CP_NUM-1:0]       cp_exception_in  // Exception signals from CPs
);

    // Coprocessor selection logic
    always_comb begin
        cp_enable = '0;
        cp_data_out = '0;
        cp_ready = 1'b0;
        cp_exception = 1'b0;
        
        if (cp_valid && cp_select < CP_NUM) begin
            cp_enable[cp_select] = 1'b1;
            cp_data_out = cp_data_from_cp[cp_select];
            cp_ready = cp_ready_in[cp_select];
            cp_exception = cp_exception_in[cp_select];
        end
    end
    
    // Forward instruction and data to selected coprocessor
    assign cp_inst_out = cp_instruction;
    assign cp_data_to_cp = cp_data_in;

endmodule

// Coprocessor MDU FSM
// Finite State Machine for Multiply/Divide Unit operations

module coprocessor_mdu_fsm #(
    parameter DATA_WIDTH = 64
)(
    input  logic                    clk,
    input  logic                    rst_n,
    
    // Control Interface
    input  logic                    mdu_start,
    input  logic [2:0]              mdu_operation,
    input  logic [1:0]              mdu_format,
    output logic                    mdu_ready,
    output logic                    mdu_busy,
    output logic                    mdu_done,
    
    // Pipeline Control
    output logic                    stage_setup_en,
    output logic                    stage_compute_en,
    output logic                    stage_normalize_en,
    output logic                    stage_complete_en,
    
    // Operation Control
    input  logic                    divide_by_zero,
    input  logic                    overflow_detected,
    output logic                    exception_raised,
    
    // Cycle Management
    output logic [4:0]              cycle_count,
    input  logic [4:0]              required_cycles,
    output logic                    operation_complete
);

    // FSM States
    typedef enum logic [2:0] {
        MDU_IDLE        = 3'b000,
        MDU_SETUP       = 3'b001,
        MDU_COMPUTE     = 3'b010,
        MDU_NORMALIZE   = 3'b011,
        MDU_COMPLETE    = 3'b100,
        MDU_EXCEPTION   = 3'b101,
        MDU_STALL       = 3'b110
    } mdu_state_t;
    
    mdu_state_t current_state, next_state;
    
    // Operation types
    typedef enum logic [2:0] {
        MDU_MUL     = 3'b000,  // Multiply
        MDU_MULH    = 3'b001,  // Multiply high
        MDU_MULHU   = 3'b010,  // Multiply high unsigned
        MDU_MULHSU  = 3'b011,  // Multiply high signed-unsigned
        MDU_DIV     = 3'b100,  // Divide
        MDU_DIVU    = 3'b101,  // Divide unsigned
        MDU_REM     = 3'b110,  // Remainder
        MDU_REMU    = 3'b111   // Remainder unsigned
    } mdu_op_t;
    
    // Internal registers
    logic [4:0]  cycle_counter;
    logic [2:0]  operation_reg;
    logic [1:0]  format_reg;
    logic        is_divide_op;
    logic        is_multiply_op;
    logic        exception_pending;
    
    // Operation classification
    always_comb begin
        is_multiply_op = (mdu_operation[2] == 1'b0); // MUL operations
        is_divide_op = (mdu_operation[2] == 1'b1);   // DIV operations
    end
    
    // State register
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            current_state <= MDU_IDLE;
            cycle_counter <= 5'b0;
            operation_reg <= 3'b0;
            format_reg <= 2'b0;
            exception_pending <= 1'b0;
        end else begin
            current_state <= next_state;
            
            // Cycle counter management
            if (current_state == MDU_COMPUTE) begin
                cycle_counter <= cycle_counter + 1;
            end else begin
                cycle_counter <= 5'b0;
            end
            
            // Latch operation parameters
            if (current_state == MDU_SETUP) begin
                operation_reg <= mdu_operation;
                format_reg <= mdu_format;
            end
            
            // Exception handling
            if ((divide_by_zero || overflow_detected) && current_state != MDU_EXCEPTION) begin
                exception_pending <= 1'b1;
            end else if (current_state == MDU_EXCEPTION) begin
                exception_pending <= 1'b0;
            end
        end
    end
    
    // Next state logic
    always_comb begin
        next_state = current_state;
        operation_complete = (cycle_counter >= required_cycles);
        
        case (current_state)
            MDU_IDLE: begin
                if (mdu_start) begin
                    next_state = MDU_SETUP;
                end
            end
            
            MDU_SETUP: begin
                if (divide_by_zero) begin
                    next_state = MDU_EXCEPTION;
                end else if (overflow_detected) begin
                    next_state = MDU_EXCEPTION;
                end else begin
                    next_state = MDU_COMPUTE;
                end
            end
            
            MDU_COMPUTE: begin
                if (exception_pending) begin
                    next_state = MDU_EXCEPTION;
                end else if (operation_complete) begin
                    next_state = MDU_NORMALIZE;
                end
                // Stay in compute state for multi-cycle operations
            end
            
            MDU_NORMALIZE: begin
                if (exception_pending) begin
                    next_state = MDU_EXCEPTION;
                end else begin
                    next_state = MDU_COMPLETE;
                end
            end
            
            MDU_COMPLETE: begin
                next_state = MDU_IDLE;
            end
            
            MDU_EXCEPTION: begin
                next_state = MDU_IDLE;
            end
            
            MDU_STALL: begin
                // Future use for pipeline stalls
                next_state = MDU_IDLE;
            end
            
            default: begin
                next_state = MDU_IDLE;
            end
        endcase
    end
    
    // Output control signals
    always_comb begin
        // Default values
        stage_setup_en = 1'b0;
        stage_compute_en = 1'b0;
        stage_normalize_en = 1'b0;
        stage_complete_en = 1'b0;
        mdu_ready = 1'b0;
        mdu_busy = 1'b0;
        mdu_done = 1'b0;
        exception_raised = 1'b0;
        
        case (current_state)
            MDU_IDLE: begin
                mdu_ready = 1'b1;
            end
            
            MDU_SETUP: begin
                stage_setup_en = 1'b1;
                mdu_busy = 1'b1;
            end
            
            MDU_COMPUTE: begin
                stage_compute_en = 1'b1;
                mdu_busy = 1'b1;
            end
            
            MDU_NORMALIZE: begin
                stage_normalize_en = 1'b1;
                mdu_busy = 1'b1;
            end
            
            MDU_COMPLETE: begin
                stage_complete_en = 1'b1;
                mdu_done = 1'b1;
            end
            
            MDU_EXCEPTION: begin
                exception_raised = 1'b1;
            end
            
            MDU_STALL: begin
                mdu_busy = 1'b1;
            end
            
            default: begin
                mdu_ready = 1'b1;
            end
        endcase
    end
    
    // Cycle count output
    assign cycle_count = cycle_counter;

endmodule

// Coprocessor MDU
// Multiply/Divide Unit for coprocessor operations

module coprocessor_mdu #(
    parameter DATA_WIDTH = 64,
    parameter ADDR_WIDTH = 64,
    parameter INST_WIDTH = 32
)(
    input  logic                    clk,
    input  logic                    rst_n,
    
    // Coprocessor Interface
    input  logic                    cp_enable,
    input  logic [INST_WIDTH-1:0]  cp_instruction,
    input  logic [DATA_WIDTH-1:0]  cp_data_in,
    output logic [DATA_WIDTH-1:0]  cp_data_out,
    output logic                    cp_ready,
    output logic                    cp_exception,
    
    // Register Interface
    input  logic [DATA_WIDTH-1:0]  rs1_data,
    input  logic [DATA_WIDTH-1:0]  rs2_data,
    output logic                    reg_write,
    output logic [4:0]              reg_addr,
    output logic [DATA_WIDTH-1:0]  reg_data,
    
    // Status and Control
    output logic [4:0]              mdu_flags,
    output logic                    mdu_busy
);

    // Instruction decode
    logic [6:0]  opcode;
    logic [4:0]  rd, rs1, rs2;
    logic [2:0]  funct3;
    logic [6:0]  funct7;
    
    assign opcode = cp_instruction[6:0];
    assign rd = cp_instruction[11:7];
    assign funct3 = cp_instruction[14:12];
    assign rs1 = cp_instruction[19:15];
    assign rs2 = cp_instruction[24:20];
    assign funct7 = cp_instruction[31:25];
    
    // MDU operation encoding
    logic [2:0] mdu_operation;
    logic [1:0] mdu_format;
    logic       mdu_start;
    logic       mdu_done;
    logic       mdu_ready_internal;
    
    // FSM interface
    logic       stage_setup_en;
    logic       stage_compute_en;
    logic       stage_normalize_en;
    logic       stage_complete_en;
    logic [4:0] cycle_count;
    logic [4:0] required_cycles;
    logic       operation_complete;
    
    // Operands and intermediate results
    logic [DATA_WIDTH-1:0]   operand_a, operand_b;
    logic [DATA_WIDTH*2-1:0] multiply_result;
    logic [DATA_WIDTH-1:0]   divide_quotient;
    logic [DATA_WIDTH-1:0]   divide_remainder;
    logic [DATA_WIDTH-1:0]   final_result;
    
    // Exception detection
    logic divide_by_zero;
    logic overflow_detected;
    logic exception_raised;
    
    // Status flags
    logic flag_zero, flag_negative, flag_overflow, flag_div_zero, flag_invalid;
    
    // Instruction decoding and operation setup
    always_comb begin
        mdu_operation = 3'b000;
        mdu_format = 2'b01; // Default 64-bit
        mdu_start = 1'b0;
        
        if (cp_enable && opcode == 7'b0110011 && funct7 == 7'b0000001) begin
            mdu_start = 1'b1;
            case (funct3)
                3'b000: mdu_operation = 3'b000; // MUL
                3'b001: mdu_operation = 3'b001; // MULH
                3'b010: mdu_operation = 3'b010; // MULHSU
                3'b011: mdu_operation = 3'b011; // MULHU
                3'b100: mdu_operation = 3'b100; // DIV
                3'b101: mdu_operation = 3'b101; // DIVU
                3'b110: mdu_operation = 3'b110; // REM
                3'b111: mdu_operation = 3'b111; // REMU
                default: mdu_start = 1'b0;
            endcase
        end else if (cp_enable && opcode == 7'b0111011 && funct7 == 7'b0000001) begin
            // 32-bit variants (RV64 *W instructions)
            mdu_start = 1'b1;
            mdu_format = 2'b00; // 32-bit
            case (funct3)
                3'b000: mdu_operation = 3'b000; // MULW
                3'b100: mdu_operation = 3'b100; // DIVW
                3'b101: mdu_operation = 3'b101; // DIVUW
                3'b110: mdu_operation = 3'b110; // REMW
                3'b111: mdu_operation = 3'b111; // REMUW
                default: mdu_start = 1'b0;
            endcase
        end
    end
    
    // Determine required cycles for operation
    always_comb begin
        case (mdu_operation)
            3'b000, 3'b001, 3'b010, 3'b011: required_cycles = 5'd3;  // Multiply operations
            3'b100, 3'b101, 3'b110, 3'b111: required_cycles = 5'd16; // Divide operations
            default:                         required_cycles = 5'd1;
        endcase
    end
    
    // Operand selection
    always_comb begin
        operand_a = rs1_data;
        operand_b = rs2_data;
    end
    
    // Exception detection
    always_comb begin
        divide_by_zero = (mdu_operation[2] == 1'b1) && (operand_b == 64'b0); // Division by zero
        overflow_detected = 1'b0;
        
        // Check for signed division overflow: -2^(n-1) / -1
        if (mdu_operation == 3'b100 || mdu_operation == 3'b110) begin // DIV or REM
            if (mdu_format == 2'b00) begin // 32-bit
                overflow_detected = (operand_a == 64'h80000000) && (operand_b == 64'hFFFFFFFF);
            end else begin // 64-bit
                overflow_detected = (operand_a == 64'h8000000000000000) && (operand_b == 64'hFFFFFFFFFFFFFFFF);
            end
        end
    end
    
    // MDU FSM instantiation
    coprocessor_mdu_fsm mdu_fsm (
        .clk(clk),
        .rst_n(rst_n),
        .mdu_start(mdu_start),
        .mdu_operation(mdu_operation),
        .mdu_format(mdu_format),
        .mdu_ready(mdu_ready_internal),
        .mdu_busy(mdu_busy),
        .mdu_done(mdu_done),
        .stage_setup_en(stage_setup_en),
        .stage_compute_en(stage_compute_en),
        .stage_normalize_en(stage_normalize_en),
        .stage_complete_en(stage_complete_en),
        .divide_by_zero(divide_by_zero),
        .overflow_detected(overflow_detected),
        .exception_raised(exception_raised),
        .cycle_count(cycle_count),
        .required_cycles(required_cycles),
        .operation_complete(operation_complete)
    );
    
    // Multiply logic
    always_comb begin
        multiply_result = 128'b0;
        case (mdu_operation)
            3'b000: begin // MUL
                if (mdu_format == 2'b00) begin // 32-bit
                    multiply_result = $signed(operand_a[31:0]) * $signed(operand_b[31:0]);
                end else begin // 64-bit
                    multiply_result = $signed(operand_a) * $signed(operand_b);
                end
            end
            3'b001: begin // MULH
                multiply_result = $signed(operand_a) * $signed(operand_b);
            end
            3'b010: begin // MULHSU
                multiply_result = $signed(operand_a) * $unsigned(operand_b);
            end
            3'b011: begin // MULHU
                multiply_result = $unsigned(operand_a) * $unsigned(operand_b);
            end
            default: multiply_result = 128'b0;
        endcase
    end
    
    // Divide logic
    always_comb begin
        divide_quotient = 64'b0;
        divide_remainder = 64'b0;
        
        if (!divide_by_zero && !overflow_detected) begin
            case (mdu_operation)
                3'b100: begin // DIV
                    if (mdu_format == 2'b00) begin // 32-bit
                        divide_quotient = {{32{1'b0}}, $signed(operand_a[31:0]) / $signed(operand_b[31:0])};
                        divide_remainder = {{32{1'b0}}, $signed(operand_a[31:0]) % $signed(operand_b[31:0])};
                    end else begin // 64-bit
                        divide_quotient = $signed(operand_a) / $signed(operand_b);
                        divide_remainder = $signed(operand_a) % $signed(operand_b);
                    end
                end
                3'b101: begin // DIVU
                    if (mdu_format == 2'b00) begin // 32-bit
                        divide_quotient = {{32{1'b0}}, operand_a[31:0] / operand_b[31:0]};
                        divide_remainder = {{32{1'b0}}, operand_a[31:0] % operand_b[31:0]};
                    end else begin // 64-bit
                        divide_quotient = operand_a / operand_b;
                        divide_remainder = operand_a % operand_b;
                    end
                end
                3'b110: begin // REM
                    if (mdu_format == 2'b00) begin // 32-bit
                        divide_remainder = {{32{1'b0}}, $signed(operand_a[31:0]) % $signed(operand_b[31:0])};
                    end else begin // 64-bit
                        divide_remainder = $signed(operand_a) % $signed(operand_b);
                    end
                end
                3'b111: begin // REMU
                    if (mdu_format == 2'b00) begin // 32-bit
                        divide_remainder = {{32{1'b0}}, operand_a[31:0] % operand_b[31:0]};
                    end else begin // 64-bit
                        divide_remainder = operand_a % operand_b;
                    end
                end
                default: begin
                    divide_quotient = 64'b0;
                    divide_remainder = 64'b0;
                end
            endcase
        end else begin
            // Handle exception cases
            if (divide_by_zero) begin
                divide_quotient = 64'hFFFFFFFFFFFFFFFF; // -1
                divide_remainder = operand_a;
            end else if (overflow_detected) begin
                divide_quotient = operand_a; // Return dividend
                divide_remainder = 64'b0;
            end
        end
    end
    
    // Result selection
    always_comb begin
        case (mdu_operation)
            3'b000: begin // MUL
                if (mdu_format == 2'b00) begin // 32-bit
                    final_result = {{32{multiply_result[31]}}, multiply_result[31:0]};
                end else begin // 64-bit
                    final_result = multiply_result[63:0];
                end
            end
            3'b001, 3'b010, 3'b011: begin // MULH variants
                final_result = multiply_result[127:64];
            end
            3'b100, 3'b101: begin // DIV, DIVU
                if (mdu_format == 2'b00) begin // 32-bit
                    final_result = {{32{divide_quotient[31]}}, divide_quotient[31:0]};
                end else begin // 64-bit
                    final_result = divide_quotient;
                end
            end
            3'b110, 3'b111: begin // REM, REMU
                if (mdu_format == 2'b00) begin // 32-bit
                    final_result = {{32{divide_remainder[31]}}, divide_remainder[31:0]};
                end else begin // 64-bit
                    final_result = divide_remainder;
                end
            end
            default: final_result = 64'b0;
        endcase
    end
    
    // Status flag generation
    always_comb begin
        flag_zero = (final_result == 64'b0);
        flag_negative = final_result[63];
        flag_overflow = overflow_detected;
        flag_div_zero = divide_by_zero;
        flag_invalid = exception_raised;
    end
    
    // Output assignments
    assign cp_data_out = final_result;
    assign cp_ready = mdu_ready_internal;
    assign cp_exception = exception_raised;
    
    assign reg_write = mdu_done && (rd != 5'b0);
    assign reg_addr = rd;
    assign reg_data = final_result;
    
    assign mdu_flags = {flag_invalid, flag_div_zero, flag_overflow, flag_negative, flag_zero};

endmodule

// Coprocessor System
// Integrates all coprocessors (CP0-CP3)
module coprocessor_system #(
    parameter ADDR_WIDTH = 64,
    parameter DATA_WIDTH = 64,
    parameter INST_WIDTH = 32,
    parameter CP_NUM = 4
)(
    input  logic                    clk,
    input  logic                    rst_n,
    
    // CPU Interface
    input  logic                    cp_valid,
    input  logic [INST_WIDTH-1:0]  cp_instruction,
    input  logic [DATA_WIDTH-1:0]  cp_data_in,
    input  logic [1:0]              cp_select,
    output logic [DATA_WIDTH-1:0]  cp_data_out,
    output logic                    cp_ready,
    output logic                    cp_exception,
    
    // System interfaces
    input  logic                    interrupt_pending,
    input  logic [DATA_WIDTH-1:0]  pc_current,
    input  logic [ADDR_WIDTH-1:0]  virtual_addr,
    input  logic [INST_WIDTH-1:0]  current_instruction,
    input  logic [ADDR_WIDTH-1:0]  mem_addr,
    input  logic [DATA_WIDTH-1:0]  mem_data,
    input  logic                    mem_write,
    input  logic                    inst_valid,
    
    // System control outputs
    output logic                    trap_enable,
    output logic [DATA_WIDTH-1:0]  trap_vector,
    output logic [ADDR_WIDTH-1:0]  physical_addr,
    output logic                    translation_valid,
    output logic                    page_fault,
    output logic                    debug_halt_request,
    output logic                    cache_flush,
    output logic                    cache_invalidate,
    
    // External interfaces
    input  logic                    external_debug_req,
    input  logic [DATA_WIDTH-1:0]  page_table_base,
    input  logic                    vm_enable,
    
    // Floating point register interface
    output logic                    fp_reg_write,
    output logic [4:0]              fp_reg_waddr,
    output logic [DATA_WIDTH-1:0]  fp_reg_wdata,
    output logic [4:0]              fp_reg_raddr1,
    output logic [4:0]              fp_reg_raddr2,
    input  logic [DATA_WIDTH-1:0]  fp_reg_rdata1,
    input  logic [DATA_WIDTH-1:0]  fp_reg_rdata2
);

    // Individual coprocessor signals
    logic [DATA_WIDTH-1:0] cp0_data_out, cp1_data_out, cp2_data_out, cp3_data_out;
    logic cp0_ready, cp1_ready, cp2_ready, cp3_ready;
    logic cp0_exception, cp1_exception, cp2_exception, cp3_exception;
    logic cp0_enable, cp1_enable, cp2_enable, cp3_enable;
    
    // System control signals from coprocessors
    logic cp0_trap_enable, cp2_debug_halt;
    logic [DATA_WIDTH-1:0] cp0_trap_vector;
    logic [ADDR_WIDTH-1:0] cp2_physical_addr;
    logic cp2_translation_valid, cp2_page_fault;
    logic cp3_cache_flush, cp3_cache_invalidate;
    
    // Coprocessor selection logic
    always_comb begin
        cp0_enable = 1'b0;
        cp1_enable = 1'b0;
        cp2_enable = 1'b0;
        cp3_enable = 1'b0;
        
        if (cp_valid) begin
            case (cp_select)
                2'b00: cp0_enable = 1'b1;  // System Control & Status (CP0)
                2'b01: cp1_enable = 1'b1;  // Floating Point Unit (CP1)
                2'b10: cp2_enable = 1'b1;  // Memory Management (CP2)
                2'b11: cp3_enable = 1'b1;  // Debug & Performance (CP3)
            endcase
        end
    end
    
    // Output multiplexing based on coprocessor selection
    always_comb begin
        case (cp_select)
            2'b00: begin
                cp_data_out = cp0_data_out;
                cp_ready = cp0_ready;
                cp_exception = cp0_exception;
            end
            2'b01: begin
                cp_data_out = cp1_data_out;
                cp_ready = cp1_ready;
                cp_exception = cp1_exception;
            end
            2'b10: begin
                cp_data_out = cp2_data_out;
                cp_ready = cp2_ready;
                cp_exception = cp2_exception;
            end
            2'b11: begin
                cp_data_out = cp3_data_out;
                cp_ready = cp3_ready;
                cp_exception = cp3_exception;
            end
            default: begin
                cp_data_out = '0;
                cp_ready = 1'b0;
                cp_exception = 1'b0;
            end
        endcase
    end
    
    // System control output assignments
    assign trap_enable = cp0_trap_enable;
    assign trap_vector = cp0_trap_vector;
    assign physical_addr = cp2_physical_addr;
    assign translation_valid = cp2_translation_valid;
    assign page_fault = cp2_page_fault;
    assign debug_halt_request = cp2_debug_halt;
    assign cache_flush = cp3_cache_flush;
    assign cache_invalidate = cp3_cache_invalidate;
    
    // CP0 - System Control and Status Register coprocessor
    coprocessor_cp0 #(
        .DATA_WIDTH(DATA_WIDTH),
        .ADDR_WIDTH(ADDR_WIDTH),
        .INST_WIDTH(INST_WIDTH)
    ) cp0_inst (
        .clk(clk),
        .rst_n(rst_n),
        .cp_enable(cp0_enable),
        .cp_instruction(cp_instruction),
        .cp_data_in(cp_data_in),
        .cp_data_out(cp0_data_out),
        .cp_ready(cp0_ready),
        .cp_exception(cp0_exception),
        .interrupt_pending(interrupt_pending),
        .pc_current(pc_current),
        .trap_enable(cp0_trap_enable),
        .trap_vector(cp0_trap_vector),
        .privilege_mode(),  // Not connected for now
        .debug_mode(),      // Not connected for now
        .debug_pc()         // Not connected for now
    );
    
    // CP1 - Floating Point Unit coprocessor
    coprocessor_cp1 #(
        .DATA_WIDTH(DATA_WIDTH),
        .ADDR_WIDTH(ADDR_WIDTH),
        .INST_WIDTH(INST_WIDTH)
    ) cp1_inst (
        .clk(clk),
        .rst_n(rst_n),
        .cp_enable(cp1_enable),
        .cp_instruction(cp_instruction),
        .cp_data_in(cp_data_in),
        .cp_data_out(cp1_data_out),
        .cp_ready(cp1_ready),
        .cp_exception(cp1_exception),
        .fp_reg_write(fp_reg_write),
        .fp_reg_waddr(fp_reg_waddr),
        .fp_reg_wdata(fp_reg_wdata),
        .fp_reg_raddr1(fp_reg_raddr1),
        .fp_reg_raddr2(fp_reg_raddr2),
        .fp_reg_rdata1(fp_reg_rdata1),
        .fp_reg_rdata2(fp_reg_rdata2),
        .fp_invalid(),      // Not connected for now
        .fp_divide_by_zero(), // Not connected for now
        .fp_overflow(),     // Not connected for now
        .fp_underflow(),    // Not connected for now
        .fp_inexact()       // Not connected for now
    );
    
    // CP2 - Memory Management Unit coprocessor
    coprocessor_cp2 #(
        .DATA_WIDTH(DATA_WIDTH),
        .ADDR_WIDTH(ADDR_WIDTH),
        .INST_WIDTH(INST_WIDTH)
    ) cp2_inst (
        .clk(clk),
        .rst_n(rst_n),
        .cp_enable(cp2_enable),
        .cp_instruction(cp_instruction),
        .cp_data_in(cp_data_in),
        .cp_data_out(cp2_data_out),
        .cp_ready(cp2_ready),
        .cp_exception(cp2_exception),
        .virtual_addr(virtual_addr),
        .physical_addr(cp2_physical_addr),
        .translation_valid(cp2_translation_valid),
        .page_fault(cp2_page_fault),
        .cache_flush(cp3_cache_flush),      // CP2 actually handles cache control
        .cache_invalidate(cp3_cache_invalidate), // CP2 actually handles cache control
        .cache_addr(),      // Not connected for now
        .page_table_base(page_table_base),
        .vm_enable(vm_enable),
        .tlb_miss(),        // Not connected for now
        .protection_fault() // Not connected for now
    );
    
    // CP3 - Debug and Performance coprocessor
    coprocessor_cp3 #(
        .DATA_WIDTH(DATA_WIDTH),
        .ADDR_WIDTH(ADDR_WIDTH),
        .INST_WIDTH(INST_WIDTH)
    ) cp3_inst (
        .clk(clk),
        .rst_n(rst_n),
        .cp_enable(cp3_enable),
        .cp_instruction(cp_instruction),
        .cp_data_in(cp_data_in),
        .cp_data_out(cp3_data_out),
        .cp_ready(cp3_ready),
        .cp_exception(cp3_exception),
        .debug_pc(pc_current),
        .debug_instruction(current_instruction),
        .debug_mem_addr(mem_addr),
        .debug_mem_data(mem_data),
        .debug_mem_write(mem_write),
        .debug_inst_valid(inst_valid),
        .debug_halt_request(cp2_debug_halt),
        .debug_single_step(), // Not connected for now
        .debug_breakpoint_hit(), // Not connected for now
        .debug_watchpoint_hit(), // Not connected for now
        .external_debug_req(external_debug_req),
        .external_halt_req(1'b0), // Not connected for now
        .debug_status(),    // Not connected for now
        .debug_halt_pc()    // Not connected for now
    );

endmodule