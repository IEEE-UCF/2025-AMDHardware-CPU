module interconnect;
endmodule
